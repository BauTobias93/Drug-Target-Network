name|status|tar|enz|tra|car
Drug1|ok|TAR1:::inh:9.5:D;TAR2:::inh:8:D;TAR3:::inh:7:D;TAR4:::inh:6:D;TAR5:::inh:8:D|||
Drug2|ok|TAR6:::inh:9.5:D;TAR7:::inh:7:D;TAR8:::inh:6:D;TAR9:::inh:8:D;TAR10:::inh:8.5:D|||
Drug3|ok|TAR1:::inh::D;TAR2:::inh::D;TAR3:::inh::D;TAR4:::inh::D;TAR5:::inh::D|||
Drug4|ok|TAR1:::inh:9.5:D;TAR2:::inh:8:D;TAR3:::inh:7:D;TAR4:::inh:6:D;TAR5:::inh:8:D|||
Drug5|ok|TAR1:::inh::D;TAR2:::inh::D;TAR3:::inh::D;TAR4:::inh:7:D|||
Drug6|ok|TAR6:::inh:5:D;TAR7:::inh:5:D;TAR8:::inh:5:D|||
Drug7|ok|TAR1:::inh:9.5:D;TAR2:::inh::D|||
Drug8|ok|TAR1:::inh:10:D;TAR2:::inh:10:D;TAR3:::inh:10:D;TAR4:::inh:10:D;TAR5:::inh:10:D;TAR6:::inh:10:D;TAR7:::inh:10:D;TAR8:::inh:10:D;TAR9:::inh:10:D;TAR10:::inh:10:D|||
Drug9|ok|TAR1:::inh::D;TAR2:::inh::D;TAR3:::inh::D;TAR4:::inh::D;TAR5:::inh::D;TAR6:::inh::D;TAR7:::inh::D;TAR8:::inh::D;TAR9:::inh::D;TAR10:::inh::D|||
