name|status|tar|enz|tra|car
Lepirudin|ok|THRB:::inh::D|||
Cetuximab|ok|EGFR:::ant::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;C1S;FCGR1;FCG2A;FCG2B;FCG2C|||
Dornase_alfa|ok|DNA|||
Denileukin_diftitox|ok_inv|IL2RA:::bin::D;IL2RB:::ago::D;IL2RG|||
Etanercept|ok_inv|TNFA:::abo::D;TNR1B;FCGR1;FCG3A;FCG2A;FCG2B;FCG2C;TNFB;FCG3B;C1S;C1R;C1QA;C1QB;C1QC|||
Bivalirudin|ok_inv|THRB:::inh::D|PERM:::inh::D||
Leuprolide|ok_inv|GNRHR:::ago:9.54:DC;GNRHR::RAT::9.3:C|CP3A4:::sub::D||
Peginterferon_alfa_2a|ok_inv|INAR2:::ago::D;INAR1:::ago::D|CP1A2:::inh::D||
Alteplase|ok|PLMN:::act::D;FIBA;UPAR;PAI1|||
Sermorelin|ok_out|GHRHR:::ago::D|||
Interferon_alfa_n1|ok_inv|INAR2:::ago::D;INAR1:::ago::D|CP1A2:::inh::D||
Darbepoetin_alfa|ok_inv|EPOR:::ago::D|||
Urokinase|ok_out|PLMN:::act::D;UPAR;UROK;TPA;PAI1;PAI2;IPSP;LRP2;ST14;NID1|||
Goserelin|ok|LSHR:::ago::D;GNRHR:::ago::D|||
Reteplase|ok_inv|PLMN:::act::D;FIBA;UPAR;PAI1|||
Erythropoietin|ok|EPOR:::ago::D|||
Salmon_Calcitonin|ok_inv|CALCR:::ago::D|||
Interferon_alfa_n3|ok_inv|INAR1:::ago::D;INAR2:::ago::D|CP1A2:::inh::D||
Pegfilgrastim|ok|CSF3R:::ago::D|ELNE:::sub::D||
Sargramostim|ok_inv|CSF2R:::ago::D;IL3RA:::ago::D;IL3RB:::ago::D;SDC2:::ago::D;PRG2|||
Peginterferon_alfa_2b|ok|INAR1:::ago::D;INAR2:::ago::D|CP1A2:::inh::D;CP2D6:::inh::D;CP2C9:::ind::D||
Asparaginase_Escherichia_coli|ok_inv|L_asparagine|||THBG:::inh::D
Thyrotropin_alfa|ok_vet|TSHR:::ago::D|||
Antihemophilic_factor_human_recombinant|ok_inv|FA10:::act::D;FA9:::cof::D;VWF:::bin::D;PAHX:::ant::D;ASGR2:::bin::D;BIP:::chap::D;CALR:::chap::D;CALX:::chap::D;LMAN1:::chap::D;LRP1:::mod::D;MCFD2:::mod::D|THRB:::act::D;PROC:::inh::D||
Anakinra|ok|IL1R1:::ant::D|||
Gramicidin_D|ok|||MDR1:::inh::D|
Human_immunoglobulin_G|ok_inv|FCGR1:::ant::D;FCGRB:::ant::D;FCG2A:::ant::D;FCG2B:::ant::D;FCG2C:::ant::D;FCG3A:::ant::D;FCG3B:::ant::D;CO3:::bin::D;CO4A:::bin::D;CO4B:::bin::D;CO5:::bin::D|||
Anistreplase|ok|PLMN:::act::D;FIBA;UPAR;PAI1|||
Insulin_human|ok_inv|INSR:::ago::D;IGF1R;RB;CBPE:::mod::D|IDE:::cli::D;NEC2:::act::D;NEC1:::act::D;CP1A2:::ind::D||
Tenecteplase|ok|PLMN:::act::D;FIBA;UPAR;PAI1;PAI2;TETN;K2C8;ANXA2;CALR;CALX;LRP1|||
Menotropins|ok|FSHR:::bin::D;LSHR|||
Interferon_gamma_1b|ok_inv|INGR1:::bin::D;INGR2:::bin::D|CP1A2:::inh::D||
Interferon_alfa_2a_Recombinant|ok_inv|INAR1;INAR2|CP1A2:::inh::D||
Desmopressin|ok|V1BR::RAT::9.7:C;V1BR::::9.43:DC;V2R::RAT::9.1:C;OXYR::RAT::9.01:C;V1AR::::8.42:DC;V2R:::ago:8.3:DC;OXYR::::8.3:C;V1AR::RAT::7.97:C|PGH2:::ind::D;PGH1:::ind::D||
Coagulation_factor_VIIa_Recombinant_Human|ok|FA10;HEPS;TFPI1;VKGC;FA7;TF|||
Oprelvekin|ok_inv|I11RA:::ago::D|||
Palifermin|ok|FGFR2:::bin::D;NRP1;FGFR1;FGFR4;FGFR3;PGBM|||
Glucagon|ok|GLR:::ago:10.15:DC;GLR::RAT::8.82:C;GLP1R:::ago:8.48:DC;GLP2R:::ago::D|||
Aldesleukin|ok|IL2RB:::ago::D;IL2RA:::ago::D;IL2RG:::ago::D|PGH2:::ind::D;PA24A:::ind::D;CP3A4:::inh::D;XDH:::ind::D;CP2E1:::inh::D||
Botulinum_Toxin_Type_B|ok_inv|VAMP2:::bin::D;VAMP1:::bin::D;SYT2|||
Omalizumab|ok_inv|FCERA:::inh::D;FCERB:::inh::D|||
Lutropin_alfa|ok|LSHR:::ago::D|||
Lyme_disease_vaccine_recombinant_OspA|ok_out|TLR2|||
Insulin_lispro|ok|INSR:::ago::D;IGF1R|CP1A2:::ind::D||
Insulin_glargine|ok|INSR:::ago::D;IGF1R|CP1A2:::ind::D||
Collagenase_clostridium_histolyticum|ok_inv|CO1A1;CO2A1;CO3A1;CO1A2|||
Rasburicase|ok_inv|Uric_acid:::met::D|||
Cetrorelix|ok_inv|GNRHR:::ant:8.9:DC;LSHR|||
Adalimumab|ok|TNFA:::abo::D|||
Somatotropin|ok_inv|GHR:::bin::D;PRLR|||
Imiglucerase|ok|Glucocerebroside|||
Abciximab|ok|ITB3:::ant::D;ITA2B:::ant::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;C1S;FCGR1;FCG2A;FCG2B;FCG2C;VTNC|||
Drotrecogin_alfa|ok_out|FA8;FA5;PAI1;TRBM;PROS;CERU;THRB;PLF4;IPSP;SPB6;VKGC;EPCR|||
Gemtuzumab_ozogamicin|ok_inv|CD33:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;C1S;FCGR1;FCG2A;FCG2B;FCG2C|||
Indium_In_111_satumomab_pendetide|exp_out|Tumor|||
Alpha_1_proteinase_inhibitor|ok|ELNE:::inh::D|||
Pegaspargase|ok_inv|L_asparagine|||THBG:::inh::D
Interferon_beta_1a|ok_inv|INAR1:::ago::D;INAR2|CP1A2:::inh::D||
Pegademase|ok|Adenosine:::met::D;GRB2:::bin::D|||
Albumin_human|ok|Nitric_oxide:::bin::D|||
Eptifibatide|ok_inv|ITB3::::6.85:DC|||
Infliximab|ok|TNFA:::inh::D|||
Follitropin|ok|FSHR:::ago::D|||
Vasopressin|ok|V2R:::ago:10.3:DC;V1AR::RAT::10.2:C;V1AR::::9.63:DC;V1BR::RAT::9.54:C;V2R::RAT::9.35:C;V1BR::::9.31:DC;OXYR::RAT::8.93:C;V2R::BOVIN::8.82:C;OXYR::::8.78:C;V2R::PIG::8.48:C||MRP2:::sub::D|
Interferon_beta_1b|ok|INAR1:::ago::D;INAR2:::ago::D|CP1A2:::inh::D||
Interferon_alfacon_1|ok_inv|INAR1:::bin::D;INAR2:::bin::D|CP1A2:::inh::D||
Hyaluronidase_ovine|ok_inv|Hyaluronan;TGFB1:::inh::D|||ALBU:::inh::D
Insulin_pork|ok|INSR:::bin::D;IGF1R;IDE;DQA2;DQB1;RB;CATD;CBPE;NEC2;NEC1;CCN3;LRP2;IBP7;SYTL4|CP1A2:::ind::D||
Trastuzumab|ok_inv|ERBB2:::abo::D;EGFR;C1R;C1QA;C1QB;C1QC;C1S;FCGR1;FCG2A;FCG2B;FCG2C;FCG3B;FCG3A|||
Rituximab|ok|CD20:::abo::D|||
Basiliximab|ok_inv|IL2RA:::abo::D;IL2RB:::abo::D;FCGR1;FCG3A;FCG2A;FCG2B;FCG2C;FCG3B;C1S;C1R;C1QA;C1QB;C1QC|||
Muromonab|ok_inv|CD3D;CD3E:::bin::D;CD3G;CD3Z;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;C1S;FCGR1;FCG2A;FCG2B;FCG2C|||
Digoxin_Immune_Fab_Ovine|ok|Digoxin|||
Ibritumomab_tiuxetan|ok_inv|CD20:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;C1S;FCGR1;FCG2A;FCG2B;FCG2C|||
Daptomycin|ok_inv|Bacterial_outer_membrane::Bacteria:destbz::D|||
Tositumomab|ok_inv|CD20:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C|||
Pegvisomant|ok|GHR:::ant::D|CP27A:::ind::D;GLNA:::inh::D;CP2CI:::inh::D;CP3A4:::ind::D;CHLE:::inh::D;CP4AB:::inh::D||
Botulinum_toxin_type_A|ok_inv|SNP25:::inh::D;RHOB|||
Pancrelipase|ok_inv|Dietary_fat:::cli::D;Dietary_protein:::cli::D;Dietary_starch:::cli::D|||
Streptokinase|ok_inv|PLMN:::act::D;PAR1:::cli::D|PA24A:::ind::D||
Alemtuzumab|ok_inv|CD52:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C|||
Alglucerase|ok_inv|Glucocerebroside|||
Capromab_pendetide|ok|FOLH1|||
Laronidase|ok|Iduronic_acid|||
Cyclosporine|ok_inv_vet|PPIA::::8.7:DC;PPID::::8.59:C;PP2BA::::8.4:C;IL2::MOUSE::8.3:C;FKB1B::::8.22:C;PPIB::::8.06:C;FKBP4::::7.8:C;FKB1A::::7.7:C;ABCBB::RAT::6.52:C;PK3CG::MOUSE::6.24:C;MDR1B::MOUSE::6.15:C;NK2R::::5.86:C;MRP2::RAT::5.71:C;CAC1C::CAVPO::5.7:C;MRP1::::5.57:C;MDR1A::MOUSE::5.44:C;PPIF:::bin::D;CANB2:::inh::D;CAMLG:::bin::D|CP3A4:::duo:6.52:DC;CP2CJ:::inh:5.15:DC;CP2D6:::inh::D;CP2C9:::inh::D;CP3A5:::inh::D;CP3A7:::ind::D|MDR1:::duo:7.7:DC;SO1B1:::inh:6.7:DC;ABCBB:::inh:6.3:DC;ABCG2:::inh:6.3:DC;NTCP:::inh:6.:DC;SO1B3:::inh:5.92:DC;MRP2:::inh:5.33:DC;MRP7:::inh::D;S22A6:::inh::D;NTCP2:::inh::D;SO1A2:::inh::D;MRP3:::inh::D|
Alefacept|ok_out|CD2:::inh::D;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C;FCG3B|||
Urofollitropin|ok_vet|FSHR:::ago::D|||
Efalizumab|ok_inv|ITAL:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C|||
Choriogonadotropin_alfa|ok|LSHR;FSHR:::bin::D|||
Antithymocyte_immunoglobulin_rabbit|ok|CD1A:::inh::D;HMR1:::ant::D;ITAL;CD86:::bin::D;FCG2B;CD4;ITB1;ITAV;ITB3|||
Filgrastim|ok|CSF3R:::sti::D;ELNE|||
Coagulation_Factor_IX_Recombinant|ok_inv|FA10:::act::D;FA11:::lig::D;FA7:::lig::D;FA8:::cof::D;THRB;LRP1;VKGC|||
Becaplermin|ok_inv|PGFRB;PGFRA;A2MG|||
Agalsidase_beta|ok_inv|Globotriaosylceramide:::lig::D|||
Octreotide|ok_inv|SSR1;SSR5;SSR2:::bin::D|PERM:::inh::D;CP3A4:::inh::D||
Interferon_alfa_2b|ok|INAR2:::bin::D;INAR1:::bin::D|CP1A2:::inh::D||
Abarelix|ok_out|GNRHR:::ant:9.1:DC|||
Oxytocin|ok_vet|OXYR:::ago:10.4:DC;OXYR::RAT::9.05:C;V2R::::8.14:C;V1AR::::8.:C;V1BR::::7.61:C;V2R::RAT::7.21:C;NEU1:::bin::D|PPCE:::sub::D||
Natalizumab|ok_inv|ITA4:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C;ICAM1|||
Enfuvirtide|ok_inv|Envelope_glycoprotein::9HIV1:::D|CP2CJ:::sub::D;CP2E1:::sub::D||
Palivizumab|ok_inv|FUS::HRSV1:::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C|||
Daclizumab|inv_out|IL2RA:::abo::D;IL2RB:::abo::D;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C|||
Bevacizumab|ok_inv|VEGFA;FCG3B;C1R;C1QA;C1QB;C1QC;FCG3A;FCGR1;FCG2A;FCG2B;FCG2C|||
Technetium_Tc_99m_arcitumomab|exp|CEAM1|||
Pyridoxal_phosphate|ok_inv_nutra|P2RX1::RAT::5.52:C;P2RX1::::5.:C;Alanine_glyoxylate_aminotransferase_homolog:::cof::D;Glutamic_acid_decarboxylase:::cof::D;SPTC3:::cof::D;SPCS:::cof::D;SRR:::cof::D;Hepatic_peroxysomal_alanine_glyoxylate_aminotransferase:::cof::D;SDSL:::cof::D;MOCOS:::cof::D;ALAT2:::cof::D;HEM0:::cof::D;GLYM:::cof::D;Glutamate:::cof::D;AT2L2:::cof::D;IGS10:::cof::D;SCLY:::cof::D;GADL1:::cof::D;KAT3:::cof::D;PDXD1:::cof::D;DDC_protein:::cof::D;Glutamate:::cof::D;5_aminolevulinate_synthase:::cof::D;Ornithine_aminotransferase_variant:::cof::D;Alpha:::cof::D;Selenocysteine_lyase_variant:::cof::D;Serine_hydroxymethyltransferase:::cof::D;Aspartate_aminotransferase:::cof::D;DDC:::cof::D;PYGM:::cof::D;PYGB:::cof::D;AATM:::cof::D;FTCD:::cof::D;PLPHP:::cof::D;BCAT2:::cof::D;BCAT1:::cof::D;CGL:::cof::D;SPTC1:::cof::D;PLPP:::cof::D;SPYA:::cof::D;HEM1:::cof::D;SERC:::cof::D;ALAT1:::cof::D;GCSP:::cof::D;KBL:::cof::D;SDHL:::cof::D;AZIN2:::cof::D;DCHS:::cof::D;CSAD:::cof::D;SPTC2:::cof::D;PYGL:::cof::D;THNS1:::cof::D;KAT1:::cof::D;ATTY:::cof::D;SGPL1:::cof::D;PNPO:::cof::D;GABT:::inh::D;AADAT:::cof::D;DCOR:::cof::D;OAT:::cof::D;AATC:::act::D;NFS1:::cof::D;GLYC:::cof::D;KYNU:::cof::D;CBS:::cof::D;DCE1:::cof::D;AGT2:::cof::D|||
Cyanocobalamin|ok_nutra|METH:::cof::D;MUTA:::cof::D;MTRR:::cof::D;MMAA:::bin::D;MMAC:::cof::D;MTHR:::cof::D|MMAB:::sub::D;COBU::SALTY:pro::D;Pancreatic_proteases::UNK:sub::D|AMNLS:::sub::D;TCO1:::sub::D;TCO2:::sub::D;IF:::sub::D;CUBN:::sub::D;LRP2;MRP1|
Ademetionine|ok_inv_nutra|PNMT::::5.32:C;AS3MT;CMTR1;COMT:::cof::D;METK1:::cof::D;CBS:::act::D;METK2:::cof::D;DCAM:::cof::D;GNMT:::cof::D|SPEE:::sub::D;CP2E1:::inh::D||
Pyruvic_acid|ok_inv_nutra|PYC;MOT3;MOT5;GABT:::inh::D;KPYM;ODPB;MOT7;KPYR;MOT6;AGT2;MOT8||SO2A1:::inh::D;MOT10:::inh::D;MOT1:::inh::DC;MOT2:::inh::DC;MOT4:::sub::DC|
Phenylalanine|ok_inv_nutra|CA2D1::MOUSE::6.01:C;TY3H:::bin::D;SYFB;SYFM;PH4H;SYFA;LAT2;ATTY||MOT10:::inh::D|
Biotin|ok_inv_nutra|IDE::::5.62:C;ACACA;PCCA;PYC;MCCA;ACACB;MCCB;SC5A6;BPL1;PCCB|CP1B1:::ind::D||
Choline|ok_nutra|SC5A7::MOUSE::5.8:C;ACHA7;PHOP1:::pro::D;PLD1:::pro::D;CHLE:::pro::D;PLD2:::pro::D;PCY1A:::pro::D;ACES:::pro::D;PCY1B:::pro::D|CHDH:::sub::D;CHKA:::sub::D;CLAT:::sub::D;CHKB:::sub::D;CEPT1:::sub::D|SC5A7:::sub::D;CTL3:::sub::D;CTL2:::sub::D;CTL4:::sub::D;CTL1:::sub::D;S22A4:::inh::D;S22A5:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|
L_Lysine|ok_nutra|SYK;CTR2;CTR3;CTR4;CTR1||S22A4:::inh::D;MOT10:::inh::D|
Arginine|inv_nutra|NFKB1::::6.6:C;ACM1::RAT::6.4:C;AGAL::::5.3:C;NOS2::::5.15:DC;CP2CJ::::5.:C;ASSY;CTR4;ARGI2;CTR1;ARLY;AZIN2;CTR3;NOS3||S22A4:::inh::D;MOT10:::inh::D;S22A5:::inh::D|
Ascorbic_acid|ok_nutra|ADA2B::::9.3:C;P4HTM;TMLH;EGLN3;PLOD1:::act::D;EGLN1;KDM5D;ALKB3;EGLN2;OGFD1;P3H3;P3H2;ALKB2;OGFD2;P3H1;P4HA1;AMD;DOPO;BODG;PLOD3;PAHX;PLOD2;XYLA::STRRU:::D;DNA;HYSA::STRPN:::D;LPH||S23A1:::::DC|
Aspartic_acid|ok_nutra|LEF::BACAN::5.9:C;NMDZ1::RAT::5.79:C;BLM::::5.45:C;FFP::BACIU::5.25:C;AL1A1::::5.05:C;ACY3;PURA1;ASGL1;SYDM;Argininosuccinate_synthetase_isoform_CRA_a;Aspartate_aminotransferase;EAA3;PURA2;PYR1;PUR6;ASPH;CMC1;SYDC;AATM;ACY1;ASSY;ASNS;ACY2;AATC;CMC2;LYSC;RNAS1||MOT10:::inh::D|
Ornithine|ok_nutra|OAZ3;GATM;OAZ2;CTR3;ORNT1;ARGI2;CTR1;CTR4;ORNT2;CTR2;OAZ1;ARGI1;OTC;OAT|||
L_Glutamine|ok_inv_nutra|BLM::::8.55:C;GLNA:::pro::D;PUR1:::pro::D;PYRG1:::ant::D|NADE:::sub::D;SYQ:::sub::D;PYR1:::sub::D;GFPT2:::sub::D;GATB:::sub::D;PUR4:::sub::D;KAT1:::sub::D;ASNS:::sub::D;GUAA:::sub::D;TGM7:::sub::D;TGM3:::sub::D;TGM4:::sub::D;TGM1:::sub::D;TGM3L:::sub::D;TGM5:::sub::D;TGM2:::sub::D;GLSL:::sub::D;GLSK:::sub::D;F13A:::sub::D|LAT2:::sub::D;AAAT:::sub::D;S38A3:::sub::D;MOT10:::inh::D|
Adenosine_phosphate|ok_inv_nutra|P2RY2::::7.07:C;SRC::::7.:C;F16P1:::ant_allo:6.85:DC;AA1R::::6.3:C;F16P1::PIG::5.89:C;P2RY1::::5.82:C;AAKG1::::5.82:C;P2RY1::MELGA::5.55:C;ADK:::pro::D;ACSL1:::pro::D;ADCY1:::pro::D;AAKB2:::act::D;AAPK1:::act::D;ACSA:::pro::D;ACS2L:::pro::D;PDE4D:::pro::D;HINT1:::pro::D;AAKB1:::act::D;PYGL:::act::D;PDE4B:::pro::D;PIM1:::pro::D;DNA;CREB1:::act::D|APT:::sub::D;AMPD1:::sub::D||
alpha_Linolenic_acid|ok_inv_nutra|NR1I2::::8.7:C;PPARA::::8.1:DC;LOX15::::6.9:C;RECQ1::::5.75:C;PPARG::::5.7:DC;FFAR4::::5.59:C;FFAR1::::5.54:C;AL1A1::::5.45:C;PGH1::::5.4:C;TYDP1::::5.3:C;AMPC::ECOLI::5.3:C;TAU::::5.05:C;RXRA;PPARD;NR1H4:::ago::D;ELOV4;TRPV1;NAC1;FADS2:::lig::D;FADS1:::lig::D|||FABP7
Methionine|ok_nutra|BHMT2:::pro::D;BHMT1:::pro::D;MAP2:::pro::D;METH:::pro::D;MTRR:::pro::D|MAT2B:::sub::D;SYMM:::sub::D;SYMC:::sub::D;MSRA:::sub::D;MSRB1:::sub::D;METK1:::sub::D;MSRB2:::sub::D;METK2:::sub::D;MTHR:::inh::D;GLNA:::inh::D|MOT10:::inh::D|
Tyrosine|ok_inv_nutra|ATTY;SYYC;SYYM;TY3H:::bin::D||MOT10:::inh::D;MOT8:::inh::D|
Calcitriol|ok_nutra|VDR:::ant:11.:DC;VDR::CHICK::10.6:C;VDR::RAT::10.4:C;VDR::BOVIN::10.3:C;VDR::PIG::10.15:C;VDRA::DANRE::8.26:C;RORG::MOUSE::5.:C;FRIL::HORSE::5.:C;HXA10|CP3A4:::sub_ind::D;CP24A:::sub_ind::D||VTDB:::bin:7.62:DC
Lutein|ok_inv_nutra||||ALBU
Cystine|ok_nutra|SLC31;BAT1;CTNS;XCT||MOT10:::inh::D|
Succinic_acid|ok_nutra|LMNA::::6.5:C;EGLN1::::5.52:C;P3H3;P3H2;P3H1;ASPH;PLOD1;SCOT1;SUCA;SSDH:::inh::D;SDHB;P4HA1;BODG;PLOD3;P4HA2;DHSD;SUCB2;S13A1;S13A2;S13A3;H17B6;SDHA;DIC;SUCB1;TMLH;SCOT2;SUCR1;C560||S22A8:::sub::D|
Riboflavin|ok_inv_nutra_vet|RBP::CHICK::8.3:C;BRCA1::::5.1:C;AL1A1::::5.05:C;IMPA1::RAT::5.:C;BLVRB:::pro::D;RISA::ECOLI:::D;RIFK:::lig::D|MTHR:::cof::D;AOFA:::cof::D|S22A6:::inh::D|
N_Acetylglucosamine|ok_inv_nutra|KLRBA::RAT::5.7:C;B4GT1;RENBP;ANAG:::act::D;NAGPA;NAGK;B4GT2;B4GT4;B4GT3|||
Glutamic_acid|ok_nutra|GRM8::::8.24:DC;GRM8::MOUSE::7.66:C;EAA3::::7.29:DC;GRM3::::7.24:C;GRM3::RAT::7.24:C;GRIK1::RAT::7.2:C;NMDZ1::RAT::7.16:C;GRIA2::RAT::6.82:C;GRIA1::RAT::6.77:C;GRM1::::6.6:DC;GRIA3::RAT::6.6:C;GRM2::::6.54:C;GRIK2::RAT::6.48:C;GRM1::RAT::6.47:C;GRIA4::RAT::6.45:C;GRM5::::6.41:C;GRIK3::RAT::6.31:C;GRM2::RAT::6.21:C;AA3R::::6.21:C;GRIK5::::6.15:DC;GRIK1::::6.15:DC;GRIK3::::6.1:DC;GRIA4::::6.06:DC;GRIA2::::6.03:DC;GRIK2::::5.96:DC;GRM7::::5.93:DC;GRM5::RAT::5.92:C;GRIA1::::5.87:DC;GRM4::::5.85:DC;GRM3:Q306L:::5.83:C;GRM2:L300Q:::5.75:C;GRM2:E273D:::5.63:C;GRM4::RAT::5.54:C;GRM8::RAT::5.47:C;GRIA3::::5.44:DC;GRM3:D279E:::5.38:C;GRM6::::5.31:C;GRM6::RAT::5.12:C;P5CS;FTCD;DCE1;DCE2;FOLH1;GSH0;DHE3;SERC;CBPQ;XCT;GRID1;DNPEP;GLSL;AASS;GHC1;GHC2;ALAT2;NMD3A;AADAT;NAGS;KAT3;NADE;LGSN;SYEM;Aspartate_aminotransferase;NMDE3;NMDE2;NMDE1;AMPE;FOLC;NMDZ1;GABT;BCAT1;GUAA;DHE4;EAA4;GSH1;EAA2;EAA1;VKGC;ALAT1;ATTY;AATC;GLNA;ASNS;SYEP;AATM;GLSK;GATB;NMD3B;GRID2;NMDE4;BCAT2;PUR4;OPLA;EAA5;GRIK4||MOT1:::sub::D;MOT10:::inh::D|
Glutathione|ok_inv_nutra|GSTK1::::7.7:DC;CP3A4;MMP9;ALDR;GPX3:::cof::D;GPX5:::cof::D;MAAI;GSTT1;GPX2:::cof::D;GPX1:::cof::D;GSTO1;GSTP1;GSTA5;GSTM4;GSTA4;GSTM3;GSTA3;GSTM1;GSHB;GSHR;LTC4S;LGUL;GLRX2;GSTO2;MGST2;GPX7:::cof::D;GPX8;Glutathione_peroxidase;GLO2;GPX6:::cof::D;GSTM5;GPX4:::cof::D;GLRX1;GSTM2;GGT1;ESTD;MGST1;TXD12;HPGDS;MGST3|GSTA2:::sub::DC;GSTA1:::sub::DC|MRP5:::sub::D;MRP4:::sub::D;MRP3:::sub::D;MRP2:::inh::D;MRP1:::inh::D|
Phosphatidyl_serine|ok_inv_nutra|DGKG;DGKD;PTSS2;NSMA3;NSMA2;AT8A1;KPCA;PTSS1;PISD;SCRB1|||
Glycine|ok_nutra_vet|NMDZ1::RAT::7.17:C;GATM;GNMT;GLRA2;GLRA3;GLYC;GLRB;SPYA;GLRA1;SC6A9;GCSP;NMD3B;SC6A5;SOX;VIAAT;AGT2;GLYL1;GLYL2;GLYM;S36A1;GLYAT;Serine_hydroxymethyltransferase;NMDE3;GSHB;GPR18;BAAT;NMDE1:::ant::D;GARS;GCSH;HEM0;HEM1;KBL||MOT10:::inh::D|
Calcifediol|ok_nutra|RORG::MOUSE::5.4:C;VDR:::ago::D|CP24A:::sub::D;CP27B:::sub::D||
Creatine|ok_inv_nutra|GAMT:::pro::D;SC6A8;KCRS:::lig::D;KCRB:::lig::D;KCRU:::lig::D;KCRM:::lig::D||S22A5:::inh::D|
Tryptophan|ok_nutra_out|MEN1::::5.15:C|I23O1:::sub::D;TPH2:::sub::D;TPH1:::sub::D;DDC:::sub::D;T23O:::sub::D;SYWC:::inh::DC;SYW::GEOSE:inh::DC;SYWM:::inh::DC|MOT10:::inh::D;MOT8:::inh::D|
Cysteine|ok_nutra|CDO1;NFS1;CSAD;SYCM;S19A3;GSHB;MGMT;SYCC;CBS;CGL;AATC;GSH1;GSH0||MOT10:::inh::D|
Thiamine|ok_inv_nutra_vet|S19A2:::bin::D;TPK1:::lig::D|CP4B1:::ind::D|S22A5:::inh::D;S22A1:::sub::D;S22A2:::inh::D|
Ergocalciferol|ok_nutra|AMPC::ECOLI::5.25:C;CCG1,CCG2,CCG3,CCG4,CCG5,CCG6,CCG7,CCG8,CA2D1,CA2D2,CA2D3,CA2D4,CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1B,CAC1A,CAC1E,CAC1G,CAC1H,CAC1I:::ind::D;VDR:::ago::D|CP11A:::sub::D;RPE:::sub::D;CP2R1:::sub::D;CP27A:::sub::D;CP27B:::sub::D;CP24A:::sub::D||VTDB:::bin::D
Citrulline|ok_inv_nutra|PADI4;PADI2;PADI3;PADI1;PADI6;NOS3;NOS2;NOS1;OTC;DDAH1;Argininosuccinate_synthetase_isoform_CRA_a;DDAH2;ASSY||S22A6:::sub::D|
Threonine|ok_nutra|SYTM;SYTC;THNS1||MOT10:::inh::D|
NADH|ok_nutra|UGDH;ADH1A;DHSO;ADH4;ADH1G;ADH1B;ADH7;GPDA;LDH6A;ADHX;ALDR;HCD2;MDHM;LDHA;MAOM;DHB4;LDH6B;LDHC;LDHB;ECHP;HCDH;MAON;BDH;MDHC;3HIDH;DHB3;HMDH;MAOX;SERA;DHB7;IDH3G;IDH3B;IDH3A;DHB1;DHB2;RDH5;G6PE;DHB8;AK1C4;IMDH2;AK1C3;PGDH;FCL;AK1C1;DHI1;3BHS2;3BHS1;IMDH1;ECHA;ALDH2;DHI2;AK1C2;NSDHL;AL3B2;MMSA;AL3A1;AL1A1;G3PT;AL9A1;AL1A3;AL1B1;AL3B1;G3P;AL1A2;AL3A2;SSDH;AL7A1;BLVRB;P5CR2;P5CR1;DHE3;ODPB;ODPAT;ODPA;BIEA;ACADS;DYR;ODO1;DHE4;DHCR7;NQO2;NU2M:::bin::D;AASS;NU3M:::bin::D;NDUS7;C1TC;MTDC;AL4A1;NB5R3;NDUAB;NU4M;DHPR;NU1M:::bin::D;NNTM;NDUA5;NDUA9;NU4LM;NDUAA;NDUA7;NDUA1;NU6M;NU5M;NDUA4;NDUA6;ACPM;NDUA2;NDUA8;NDUA3;NDUB8;NDUC2;NDUB1;NDUS1;NDUBA;NDUB4;NDUB3;NDUB2;NDUB7;NDUB9;NDUS2;NDUB5;NDUC1;NDUB6;NDUV3;DLDH;NDUS3;GSHR;NDUAC;NDUS5;NDUS4;NDUV1;NDUV2;NDUAD;CDO1;NDUS6;NUA4L;NDUS8;CP4AB;ODP2;GCST;MSMO1;HMOX1;HMOX2;CP17A;TYRO|XDH:::sub::D;AOXA:::sub::D;ADH6:::act::D;AK1A1:::sub::D;ADH1A:::sub::D;ADH1B:::sub::D;ADH4:::sub::D;ADHX:::sub::D;ADH7:::sub::D||
Folic_acid|ok_nutra_vet|TSHR::::5.1:C;KDM4E::::5.:C;FOLR1;FOLR2:::bin::D;FOLR3:::bin::D|DYR:::sub::D;MTHR:::sub::D;GGH:::sub::D|MFTC:::sub::D;PCFT:::sub::D;ABCG2:::sub::D;MRP4:::inh::D;S22A6:::inh::D;MRP3:::sub::D;ABCCB:::sub::D|
Icosapent|ok_nutra|PPARA::::5.96:DC;PPARG:::ago:5.8:DC;OXER1::::5.7:C;PPARD:::ago:5.4:DC;PGH2::SHEEP::5.15:C;TRPV1:::ind::D;NAC1:::inh::D;FFAR1:::ago::D;ACSL3:::ind::D;ACSL4:::ind::D;FADS1:::ago::D;PGH1:::inh::D;PGH2:::inh::D|||ALBU;FABP7:::ago::D
Valine|ok_nutra||SYVC:::sub::DC;BCAT1:::sub::DC;PCCB:::sub::DC|MOT10:::inh::D|
Vitamin_A|ok_nutra_vet|LACB::BOVIN::7.44:C;AL1A1::::5.22:DC;HPGDS;APOD;RLBP1;AL1A2;RET3;RDH13;RDH5;RET1;LRAT;RDH8;RDH14;DHRS4;RDH11;RETST;AL1A3;DHRS3;RDH12|CP26A:::sub_ind::D||RET4::::6.74:DC;ALBU;RET2;RET7;RET5
Vitamin_E|ok_nutra_vet|LMNA::::6.95:C;TAU::::5.45:C;S14L4;PP2AA;PP2AB;DGKA;KPCA;LOX5;KPCB;NR1I2|CP3A4:::sub_ind::D;SODC:::ind::D;HMOX1:::ind::D;NQO1:::ind::D;GSH1:::ind::D;GSTM3:::ind::D;GSTO1:::inh::D;GSTP1:::inh::D;GSTA2:::ind::D|ABCG1;NPCL1;ABCA1:::tra::D;SCRB1:::tra::D|TTPA::::5.62:DC;PLTP:::car::D;S14L2:::car::DC;S14L3:::car::DC
Pyridoxine|ok_inv_nutra_vet|PDXK:::lig::D|CP1A1:::inh::D||
Lipoic_acid|ok_inv_nutra|ACES::::9.:C;LMNA::::6.45:C;THB::::6.05:C;END4::ECOLI::6.05:C;NR1I2::::5.55:C;BLM::::5.1:C;SC5A6;LIAS;LIPT|NCPR:::inh::D||
Cholecalciferol|ok_nutra|VDR:::ago:9.68:DC;GLRA1::::6.4:C;RORG::MOUSE::5.35:C|CP2C8:::inh::D;CP1A1:::inh::D;CP11A:::sub::D;CP3A4:::sub::D;CP2J2:::sub::D;CP27A:::sub::D;CP2R1:::sub::D||VTDB
Menadione|ok_nutra|AOXA::MACFA::6.96:C;AOXA::MOUSE::6.82:C;AOXA::RAT::6.72:C;AOFB::::6.4:C;I23O1::::6.:C;AOXA::RABIT::5.7:C;MPIP2::::5.66:C;CP2CJ::::5.6:C;TAU::::5.3:C;AMPC::ECOLI::5.25:C;CP2C9::::5.2:C;ALDOA::RABIT::5.2:C;RORG::MOUSE::5.2:C;UBP2::::5.2:C;CP2D6::::5.1:C;ABHD5::::5.1:C;PLIN5::::5.02:C;P53::::5.:C;G3P::::5.:C;OSTCN:::ago::D;NQO1;NQO2;PROZ:::act::D;PROS:::act::D;PROC:::act::D;FA10:::act::D;FA9:::act::D;FA7:::act::D;THRB:::act::D;VKORL:::cof::D;VKOR1:::cof::D;VKGC:::cof::D|CP1A2:::ind:6.8:DC;AOXA:::inh:6.7:DC;CP2A6:::inh::D;CP1A1:::duo::D;MTHR:::sub::D;XDH:::sub::D||
Adenine|ok_nutra|LMNA::::5.6:C;COBT::SALTY:::D;MTAP;DNA;RUVB::THET8:::D;SRPK2;Nucleoside_2_deoxyribosyltransferase::LACHE:::D;MUTY::ECOLI:::D;PECR;PPAC;ACACB;MTNN::ECOLI:::D;APT|UD11:::inh::D||
Asparagine|ok_inv_nutra|SYNC;ASNS;S38A3;SYNM;ASGL1;AAAT||MOT10:::inh::D|
Pravastatin|ok|HMDH:::inh:8.25:DC;HMDH::RAT::7.89:C;HDAC2:::inh::D||SO1B1:::sub:5.47:DC;SO1B3:::sub::D;ABCBB:::sub::D;MOT1:::sub::D;S22A7:::sub::D;ABCG2:::sub::D;S22AB:::sub::D;MRP2:::sub::D;S22A8:::inh::D;S22A6:::inh::D;SO1A2:::sub::D;MDR1:::sub::D;SO2B1:::sub::D|
Fluvoxamine|ok_inv|SC6A3::::8.84:C;SGMR1::::7.44:C;SGMR1::RAT::7.44:C;SC6A4::RAT::6.27:C;KCNH2::::5.51:DC;CAC1C::CAVPO::5.31:C;IMPA1::RAT::5.:C;SC6A4:::inh::D|CP2D6:::inh:5.1:DC;CP2C9:::inh:5.07:DC;CP2B6:::inh::D;CP2CJ:::inh::D;CP3A4,CP343,CP3A5,CP3A7:::inh::D;CP3A4:::inh::D;CP1A1:::inh::D;CP1A2:::inh::D|ABCBB:::sub::D;MDR1:::inh::D|
Valsartan|ok_inv|AGTRB::RAT::8.72:C;AGTR1:::ant:8.57:DC;AGTRA::RAT::8.47:C|CP2C9:::sub::D|MRP2:::sub::D;SO1B1:::inh::D;SO1B3:::sub::D|
Ramipril|ok|ACE:::inh:8.4:DC;ACE::RABIT::6.6:C;BKRB1|CHLE:::inh::D|S15A2:::sub::D;S15A1:::sub::D|
Masoprocol|ok_inv|SHBG|LOX5:::inh::DC||
Flunisolide|ok_inv|GCR:::ago:8.62:DC|CP3A4:::sub_ind::D||CBG:::ago::D
Baclofen|ok|GABR1::RAT::7.52:C;GBRP::RAT::7.52:C;CP3A4::::7.5:C;GABR1:::ago:7.46:DC;AA3R::::7.3:C;BLM::::6.7:C;NFKB1::::5.25:C;LMNA::::5.2:C;GABR2:::ago::D|||
Amphetamine|ok_ill_inv|SC6A3::RAT::6.02:C;SC6A2::MOUSE::6.:C;CP2A5::MOUSE::5.55:C;5HT3A::RAT::5.27:C;5HT2B::RAT::5.27:C;5HT1B::RAT::5.12:C;Vesicle_monoamine_transporter_type_2;AOFA,AOFB:::inh::D;SC6A4:::bin::D;AOFB:::inh::D;DRD2:::bin::D;ADRB1,ADRB2,ADRB3:::ago::D;ADA1A,ADA1B,ADA1D,ADA2A,ADA2B,ADA2C:::ago::D;SC6A2:::sti::D;TAAR1:::ago::D;CART:::ago::D;SC6A3:::neg::D;VMAT2:::inh::D|CP2A6:::inh:5.46:DC;CP2D6:::sub::D|S22A5:::sub::D;S22A3:::sub::D|
Pentagastrin|ok|GASR::MOUSE::9.1:C;GASR::RAT::8.17:C;GASR:::ago:7.84:DC;CCKAR::RAT::6.22:C|CHLE:::ind::D||
Nicotine|ok|ACHA3::RAT::11.:C;ACHB2:::ago:9.22:DC;ACHA4::RAT::9.08:C;ACHA::TETCF::9.:C;ACHA7:::ago:8.97:DC;ACHB2::MOUSE::8.92:C;ACHA4::CHICK::8.72:C;ACHA9::RAT::8.62:C;ACHB3::RAT::8.48:C;ACHA2::RAT::8.26:C;ACHA4::MOUSE::8.15:C;ACHA7::RAT::7.8:C;ACHB4:::ago:7.64:DC;ACHA3:::ago:7.35:DC;ACHP::LYMST::7.2:C;ACHB4::RAT::7.14:C;ACHB4::MOUSE::6.78:C;ACHA7::MOUSE::6.61:C;ACHA::::5.83:C;ACH4::DROME::5.57:C;CRTY::PANAN::5.32:C;CLAT:::inh::D;CP19A:::inh::D;ACHB3:::ago::D;ACH10:::ago::D;ACHA9:::ago::D;ACHA6:::ago::D;ACHA5:::ago::D;ACHA2:::ago::D;ACHA4:::ago::D|CP2A6:::inh:5.36:DC;AOFB:::inh::D;AOFA:::inh::D;CP3A4:::sub::D;CP2D6:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1A2:::sub_ind::D;CP1A1:::sub_ind::D;CP2B6:::sub::D;CP2AD:::sub::D;CP2E1:::duo::D|S22A4:::inh::D;S22A5:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|
Cevimeline|ok|ACM3:::ago::D;ACM1:::ago::D|CP2D6:::sub::D;CP3A4:::sub::D;FMO1:::sub::D||
Lorazepam|ok|TSPO;GABAR:::aga::D|CP3A4:::sub::D;UDB15:::sub::D||
Esmolol|ok|ADRB1:::ant:6.94:DC;ADRB2::CAVPO::5.2:C|CP2D6:::sub::D||
Bortezomib|ok_inv|PSB5:::inh:9.26:DC;PSMD1::::8.59:C;PSB8::::8.09:C;NFKB2::::8.01:C;PSB8::MOUSE::7.77:C;PSB1:::inh:7.28:DC;CTRB1::::6.49:C;CATG::::6.28:C;PSB2::::6.23:C;CAH2::::5.94:C;CMA1::::5.92:C;CAH1::::5.89:C;ELNE::::5.64:C;CTRA::BOVIN::5.62:C;PPGB::::5.04:C|CP2C9:::inh::D;CP1A2:::inh::D;CP2D6:::sub::D;CP2CJ:::inh::D;CP3A4:::sub::D||
Ethchlorvynol|ok_ill_out|GABAR:::aga::D|||
Carbidopa|ok|MK01::::7.4:C;HCD2::::6.8:C;TYDP1::::5.95:C;KDM4E::::5.65:C;LOX15::::5.4:C;AL1A1::::5.15:C;CP1A2::::5.1:C;DDC:::inh::D|||
Phentermine|ok_ill|TAAR1::::5.26:C;NPY:::inh::D;AOFB:::ant::D;AOFA:::ant::D;SC6A3:::inh::D;SC6A4:::inh::D;SC6A2:::inh::D|CP3A4:::sub::D||
Indecainide|ok|SCN5A:::inh::D|||
Tramadol|ok_inv|OPRM:::ago:6.:DC;SC6A4:::inh:5.96:DC;SC6A2:::inh:5.7:DC;ADA2A,ADA2B,ADA2C:::sti::D;AA1R:::sti::D;NMDA:::inh::D;TRPV1:::ago::D;SCN2A:::inh::D;NK1R:::inh::D;ACM1:::ant::D;ACM3:::ant::D;Alpha_7_nicotinic_cholinergic_receptor_subunit:::ant::D;OPRD:::ago::D;OPRK:::ago::D;5HT2C:::ant::D|UD11:::sub::D;CP2B6:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D|MDR1:::sub::D|
Vidarabine|ok_inv|DPP4::::7.21:C;KITH::HHV1:ind::D;KITH::VZVD:ind::D;DNA:::destbz::D;DPOL::EBVB9:inh::D|ADA:::sub::D||
Betaxolol|ok_inv|ADRB1:::ant:8.8:DC;ADRB1::RAT::8.53:C;ADRB2::CAVPO::6.98:C;ADRB2::BOVIN::6.18:C;ADRB2:::ant::D|CP2D6:::sub::D;CP1A2:::sub::D||
Fluconazole|ok_inv|CP51::MYCTU::6.7:C;LMNA::::6.3:C;HS90A::::5.33:C;CP121::MYCTU::5.22:C;CP51::CANAL:inh::D|CP3A4:::inh:5.1:DC;CP2CJ:::inh:5.09:DC;CP2C9:::inh:5.04:DC;CP3A5:::inh::D|MDR1:::inh::D|
Troglitazone|ok_out|PPARG:::ago:6.52:DC;PPARG::MOUSE::6.11:C;CAC1C::CAVPO::6.1:C;5HT2B::::6.08:C;CAH2::::6.01:C;MK01::::5.91:C;ALDR::RAT::5.69:C;AOFB::::5.68:C;THAS::::5.53:C;AA3R::::5.53:C;ABCBB::RAT::5.41:C;I23O2::MOUSE::5.35:C;AOFA::RAT::5.32:C;NR1I2::::5.16:C;CAC1C::RAT::5.02:C;GSTP1;PPARA;PPARD;ERR1:::ANT::D;ERR3:::ANT::D;S29A1:::inh::D;PAI1:::ant::D;ACSL4:::inh::D|CP2C9:::inh:5.4:DC;UDB15:::sub::D;UD2B7:::sub::D;UD110:::sub::D;UD19:::sub::D;UD18:::sub::D;UD17:::sub::D;UD16:::inh::D;UD14:::sub::D;UD13:::sub::D;CP3A7:::inh::D;CP3A5:::inh::D;CP2B6:::ind::D;CP1A1:::ind::D;CP19A:::inh::D;CP2CJ:::inh::D;UD11:::sub::D;CP2C8:::inh::D;CP3A4:::ind::D|ABCBB:::inh:5.57:DC;SO1B1:::inh::D|
Oseltamivir|ok|NRAM::INBLE::8.96:C;NRAM::I77AB::8.86:C;NRAM::I68A0::8.81:C;NRAM::I34A1::8.15:C;NEUR2:::inh::D;NEUR1:::inh::D;NRAM::I83A1:inh::D|EST1:::sub::D|S22A8:::sub::D;S15A1:::sub::D;MRP4:::sub::D|
Erythromycin|ok_inv_vet|KCNH2:::inh:7.41:DC;MTLR:::ago:7.36:DC;AMPC::ECOLI::5.7:C;23S_ribosomal_RNA::Gut_flora:inh::D|CP3A4:::inh:6.72:DC;CP3A5:::inh::D;CP3A7:::inh::D|SO1A2:::inh::D;MRP2:::sub::D;SO1B1:::inh::D;MDR1:::inh::D;ABCBB:::inh::D;SO1B3:::inh::D|
Hydroxocobalamin|ok|METH:::cof::D;MUTA:::cof::D;MTRR;MMAA;TCO1;AMNLS;CUBN;MMAB;MMAC|||TCO2:::sub::D
Caffeine|ok|ACM1::RAT::7.45:C;LEF::BACAN::6.:C;AA2AR:::ant:5.61:DC;KCNH2::::5.31:C;ACES::::5.14:C;AA2AR::RAT::5.03:C;PDE1B,PDE4D,PDE3B,PDE5A:::inh::D;AA3R:::ant::D;AA2BR:::ant::D;ATM:::inh::D;ITPR1,ITPR2,ITPR3:::inh::D;PK3CB:::inh::D;PK3CA:::inh::D;PK3CD:::inh::D;PRKDC:::inh::D;PDE1A,PDE1B,PDE1C,PDE10,PDE4A,PDE4B,PDE4C,PDE4D,PDE7B,PDE2A,PDE3A,PDE3B,PDE5A,PDE6C,PDE11,PDE7A,PDE8A,PDE8B,PDE9A,PDE6A,PDE6B:::inh::D;RYR1;PDE4B:::inh::D;AA1R:::ant::D|CP2D6:::sub::D;CP1B1:::sub::D;CP1A1:::inh::D;CP2C9:::sub::D;CP2C8:::sub::D;CP2E1:::sub::D;CP3A4:::sub::D;CP1A2:::inh::D|ABCG2:::inh::D|
Succinylcholine|ok|ACM3:::ago::D;ACM2:::ago::D;ACM1:::ago::D;Alpha_7_nicotinic_cholinergic_receptor_subunit:::ago::D;ACH10:::ago::D|CHLE:::sub::D||
Sildenafil|ok_inv|PDE5A::RAT::9.52:C;CNCG:::inh:9.3:DC;PDE5A::CANLF::9.:C;PDE5A:::inh:8.8:DC;PDE5A::BOVIN::8.22:C;PDE6B::BOVIN::7.7:C;PDE6C::::7.62:C;PDE6C::BOVIN::7.48:C;AA2AR::::6.85:C;PDE6A::BOVIN::6.85:C;PDE1C::RAT::6.59:C;PDE1A::::6.57:C;PDE1B::BOVIN::6.4:C;ADA1B::RAT::6.09:C;AA1R::::6.06:C;PDE11::::5.64:C;PDE10::::5.51:C;KCNH2::::5.48:C;PDE9A::::5.47:C;I23O2::MOUSE::5.35:C;PDE4D::RAT::5.34:C;PDE7A::::5.33:C;PDE4A::::5.3:C;PDE3A::::5.15:C;CNRG:::inh::D|CP3A4:::sub:5.3:DC;CP2E1:::inh::D;CP2D6:::sub::D;CP2CJ:::inh::D;CP2C9:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D|MRP5:::inh:5.92:DC;MDR1:::inh::D;SO1B1:::inh::D;MRP7:::inh::D;MRP4:::inh::D|
Dofetilide|ok_inv|KCNH2:::inh:8.39:DC;KCJ12:::inh::D;KCNK2:::inh::D|CP3A4:::sub::D|S22A2:::sub::D|
Pyrimethamine|ok_inv_vet|DRTS::PLAFK:inh:9.72:DC;DYR:::inh:8.1:DC;DYR::PNECA::8.01:C;DRTS:S108N:PLAFK:inh:7.54:DC;DRTS::TOXGO::7.1:C;S47A1::MOUSE::6.84:C;DYR::RAT::5.85:C;HEXB::::5.51:DC;S22A1::MOUSE::5.44:C;STRP::STRP1::5.4:C;DYR::CANAX::5.3:C;CP3A4::::5.3:C;P53::::5.1:C;CP2D6::::5.1:C;HEXA:G269S:::5.07:C;CP1A2::::5.:C|CP2C8:::inh::D|S47A2:::inh::D;S47A1:::inh::D|
Reserpine|ok_inv|VMAT2::BOVIN::9.:C;SCN1A::::5.8:C;OPRM::::5.77:C;CP3A4::::5.4:C;MDR1A::MOUSE::5.39:C;ACM1::RAT::5.25:C;END4::ECOLI::5.2:C;NORA::STAAU::5.15:C;MK01::::5.1:C;CASP7::::5.1:C;CASP1::::5.1:C;NORA:A116E:STAAU::5.04:C;NPSR1::::5.:C;BIRC5;VMAT1:::inh::D;VMAT2:::inh::D|CP3A5:::ind::D|MDR1:::duo:7.:DC;SO2B1:::inh::D;SO1B1:::inh::D;S22A2:::sub::D;MRP2:::inh::D;ABCBB:::inh::D;S22A1:::inh::D|
Azithromycin|ok|LMNA::::6.2:C;TSHR::::5.1:C;PADI4:::inh::D;23S_ribosomal_RNA::Gut_flora:inh::D|CP3A4:::inh::D|MRP2:::inh::D;MDR1:::inh::D|
Ticlopidine|ok|ADA2B::::6.86:C;ADA2A::::6.84:C;ADA2C::::6.77:C;SGMR1::::6.75:C;LMNA::::5.:C;P2Y12:::ant::D|CP2CJ:::inh:7.4:DC;CP2B6:::inh:6.7:DC;CP2D6:::inh:6.4:DC;CP1A2:::inh:6.3:DC;CP2E1:::inh::D;CP2C8:::inh::D;CP2C9:::inh::D;PERM:::sub::D||
Trospium|ok|ACM1:::ant::D|CP2D6:::inh::D||
Adapalene|ok|RARB:::ago:7.47:DC;RARG:::ago:6.89:DC;RARA:::ago:5.96:DC;GLRA1::::5.89:C;LMNA::::5.5:C;PGH2:::inh::D;RXRA;RXRB:::ago::D;RXRG:::ago::D|||
Midodrine|ok|ADA1A:::ago::D;ADA1B:::ago::D;ADA1D:::ago::D|CP2D6:::sub::D|S15A1|
Remikiren|exp|RENI:::inh:10.6:DC|||
Pantoprazole|ok|ATP4A:::inh:6.:DC;LMNA::::5.9:C;S22A2::::5.82:C;S47A1::::5.55:C;FAS::::5.39:C;DDAH1:::inh::D|CP3A4:::sub::D;CP2CJ:::inh::D|ABCG2:::inh:5.:DC;S22A8:::inh::D;MDR1:::inh::D|
Torasemide|ok|CP3A4::::6.:C;HIF1A::::5.4:C;S12A2:::inh::D;S12A1:::inh::D|CP2C9:::inh::D;CP2C8:::sub::D|SO1B1:::sub::D|ALBU:::sub::D
Citalopram|ok|SC6A4:::inh:9.32:DC;SC6A4::RAT::8.82:C;SC6A3::MOUSE::8.54:C;KCNH2::::8.:C;5HT2C::::6.81:C;SGMR1::::6.78:C;HRH1:::bin:6.43:DC;ADA1A::RAT::6.15:C;5HT2B::::5.93:C;ADA1D::::5.79:C;ADA1B::RAT::5.74:C;SC6A2::::5.66:C;SC6A3::RAT::5.03:C|CP1A2:::inh::D;CP2D6:::inh::D;CP2CJ:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Eletriptan|ok_inv|5HT7R:::ago::D;5HT2B:::ago::D;5HT1E:::ago::D;5HT1A:::ago::D;5HT1F:::ago::D;5HT1B:::ago::D;5HT1D:::ago::D|CP2A6:::ind::D;PGH1:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D|MDR1:::sub::D|
Bethanidine|ok|ADA2A:::ago::D;KCNJ1:::inh::D;ADRB1:::ant::D|||
Moxifloxacin|ok_inv|GYRB::ECOLI::6.52:C;PARC::STAAU::6.1:C;GYRB::STAAU::5.11:C;GYRA::MYCTU::5.04:C;TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A2:::inh::D||
Oxyphenonium|ok|ACM1:::ant::D|||
Nelfinavir|ok|MDR1A::MOUSE::5.64:C;OPRM::::5.23:C;DRD1::::5.19:C;FYN::::5.1:C;AA3R::::5.08:C;SC6A2::::5.06:C;NK2R::::5.01:C;HIV::9PLVG:inh::D|CP3A4:::inh:6.32:DC;CP3A5:::inh:6.24:DC;CP2D6:::inh::D;CP2C9:::inh::D;UD11:::ind::D;CP2CJ:::sub_ind::D;CP2B6:::inh::D;CP3A7:::inh::D|MDR1:::duo:6.46:DC;ABCBB:::sub::D;SO2B1:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;SO1A2:::inh::D;S22A1:::inh::D|ALBU
Isoetharine|ok|ADRB2:::ago:6.:DC;ADRB1:::ago::D|||
Glimepiride|ok|RORG::MOUSE::5.:C;ABCC8:::ind::D;KCNJ1:::inh::D;KCJ11:::inh::D|CP2C9:::sub::D|ABCBB:::sub::D|
Diflorasone|ok|GCR:::ago::D|||
Indinavir|ok|NK2R::::5.77:C;S47A1::::5.77:C;THAS::::5.73:C;S47A2::::5.11:C;Pol_polyprotein::9HIV1:inh::D|CP3A4:::inh:6.82:DC;UD11:::inh::D;CP2D6:::inh::D;CP3A5:::inh::D;CP3A7:::inh::D|ABCBB:::sub::D;SO2B1:::inh::D;MRP2:::sub::D;SO1B1:::inh::D;SO1A2:::inh::D;MRP1:::inh::D;S22A1:::inh::D;MDR1:::duo::D|
Gadodiamide|ok_inv||||
Guanadrel|ok|SC6A2:::pag::D|||
Lovastatin|ok_inv|HMDH:::inh:9.22:DC;HMDH::RAT::8.52:C;HMDH::MOUSE::7.57:C;CHLE::HORSE::5.96:C;ACES::ELEEL::5.57:C;ITAL:::inh_allo:5.42:DC;LMNA::::5.25:C;RORG::MOUSE::5.15:C;SC6A3::::5.1:C;SC6A2::::5.06:C;NK2R::::5.03:C;HIF1A::::5.:C;HDAC2|CP3A4:::inh:5.:DC;CP2CJ:::sub::D;UD2B7:::sub::D;UD13:::sub::D;UD11:::sub::D;CP2C8:::sub::D;PON3:::sub::D|MDR1:::inh:5.:DC;SO1B3;SO2B1;ABCBB:::sub::D;MRP2:::sub::D;SO1B1:::inh::D;SO1A2:::inh::D|ALBU:::sub::D
Enflurane|ok_inv_vet|ATPD;GRIA1:::ant::D;AT2C1:::inh::D;KCNA1:::ind::D;KCNN4:::inh::D;GLRA1,GLRB:::ago::D;GABAR:::aga::D|CP2E1:::sub::D||ALBU
Cefotiam|ok_inv|PBPA::CLOPE:ind::D||S22A8:::inh::D;S22A6:::inh::D|
Pregabalin|ok_inv|CA2D1||LAT1;EAA3|
Temazepam|ok_inv|LMNA::::6.55:C;GABAR:::aga::D;TSPO;GBRT:::pot::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2C9:::sub::D;CP2B6:::sub::D;CP3A4:::sub::D||
Methyclothiazide|ok|CAH4:::inh::D;CAH2:::inh::D;CAH1:::inh::D;S12A1:::inh::D|||
Aminosalicylic_acid|ok|HPPK::MYCTU:::D;PA2GE;LOX5:::inh::D;IKKA:::inh::D;PGH2:::inh::D|PERM:::inh::D||
Reboxetine|ok_exp|SC6A2:::inh::D|CP3A4:::inh::D;CP2D6:::inh::D|MDR1:::inh::D|
Milrinone|ok|BLM::::7.65:C;PDE3A:::inh:6.82:DC;PDE3B::::6.55:C;AMPC::ECOLI::6.2:C;PDE5A::::6.13:C;PDE4A::::5.96:C;TSHR::::5.4:C;PGH1::::5.33:C;PDE4A::CAVPO::5.33:C;PDE5A::BOVIN::5.3:C|||
Pipobroman|ok|CP3A4::::7.2:C;LMNA::::6.3:C;AL1A1::::6.05:C;CYSP::TRYCR::5.2:C;TYDP1::::5.1:C;MEN1::::5.:C;DNA:::cov::D|||
Butabarbital|ok_ill|GABAR:::aga::D;ACHA4:::ant::D;ACHA7:::ant::D;GRIA2:::ant::D;GRIK2:::ant::D|||
Nevirapine|ok|LMNA::::7.45:C;MK01::::5.45:C;Reverse_transcriptase_RNaseH::9HIV1:inh::D|CP3A7:::sub::D;CP1A2:::inh::D;CP2D6:::inh::D;CP2A6:::sub::D;CP2C9:::ind::D;CP3A5:::sub::D;CP3A4:::sub_ind::D;CP2B6:::sub_ind::D|S22A1:::inh::D|ALBU
Oxiconazole|ok|AA3R::::6.45:C;SC6A4::::6.37:C;ADA2C::::6.22:C;THAS::::6.21:C;DRD3::::6.17:C;ACM3::::6.02:C;CP2D6::::6.:C;NK2R::::5.97:C;ACM1::::5.94:C;5HT2A::::5.92:C;ADA2A::::5.82:C;ADA2B::::5.78:C;OPRD::::5.73:C;SC6A2::::5.72:C;SC6A3::::5.68:C;DRD1::::5.68:C;5HT2B::::5.53:C;CP2C9::::5.52:C;5HT1A::RAT::5.5:C;ADRB3::::5.45:C;ACES::::5.33:C;NR1I2:::pag::D;ERG7::CANAL:inh::D;CP51::CANAL:inh::D|CP2CJ:::sub:7.4:DC;CP3A4:::ind:7.05:DC||
Alclometasone|ok|GCR:::ago::D|CP3A4:::sub::D||CBG:::bin::D
Butalbital|ok_ill|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA4:::pot::D;GBRA5:::pot::D;GBRA6:::pot::D;ACHA4:::ant::D;ACHA7:::ant::D;GRIA2:::ant::D;GRIK2:::ant::D;GABAR:::aga::D|||
Cladribine|ok_inv|LMNA::::7.3:C;HD::::5.35:C;AA1R::RAT::5.14:C;PNPH:::ind::D;DPOE4:::inh::D;DPOE3:::inh::D;DPOE2:::inh::D;DPOE1:::inh::D;DPOLA:::inh::D;DNA;RIR2B:::inh::D;RIR2:::inh::D;RIR1:::inh::D|DCK:::sub::D|S28A3;ABCG2:::sub::D|
Ranolazine|ok_inv|SCN5A::::5.17:C;Fatty_acid::UNK:::D;ADRB1:::ant::D;ADA1A,ADA1B,ADA1D:::ant::D;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4:::inh::D;KCJ12,KCJ14,KCNJ2,KCNJ4:::inh::D;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A,SCN1B,SCN2B,SCN3B,SCN4B:::inh:,,,,,,5.17,,,,,,,:DC|CP2D6:::inh::D;CP3A4:::inh::D|MDR1:::inh::D;ABCBB:::sub::D|A1AG1:::bin::D;ALBU:::bin::D
Mesalazine|ok|TYDP1::::6.:C;RECQ1::::5.4:C;KDM4E::::5.4:C;CP2CJ::::5.3:C;CASP1::::5.2:C;CASP7::::5.1:C;CP3A4::::5.1:C;AL1A1::::5.05:C;HCD2::::5.:C;HIF1A::::5.:C;NAT::MYCTU:::D;PERM;IKKB:::inh::D;IKKA:::inh::D;PPARG:::ago::D;LOX5:::inh::D;PGH1:::inh::D;PGH2:::inh::D|ARY1:::sub::D||
Benzatropine|ok|ACM1:::ant:9.88:DC;ACM3::::9.57:C;ACM4::::9.48:C;HRH1:::ant:9.43:DC;ACM1::RAT::9.23:C;ACM5::::8.84:C;ACM2::RAT::8.59:C;ACM2::::8.44:C;5HT2A::::8.16:C;SC6A3::RAT::8.1:C;ADA1D::::7.59:C;ADA2B::::7.52:C;5HT2C::::7.49:C;ADA1B::RAT::7.39:C;ADA1A::RAT::7.24:C;ADA2C::::7.24:C;SGMR1::::7.23:C;5HT2B::::6.9:C;SC6A3:::inh:6.71:DC;ADA2A::::6.69:C;DRD3::::6.65:C;HRH2::::5.93:C;5HT6R::::5.89:C;SC6A2:::inh:5.86:DC;SC6A4::RAT::5.29:C;SC6A4:::inh::D|||ALBU:::bin::D
Ziprasidone|ok|5HT2A:::ant:10.1:DC;5HT2A::RAT::9.38:C;DRD2::RAT::9.38:C;ADA1A::RAT::9.3:C;5HT2C:::ant:9.26:DC;5HT1A:::ago:8.8:DC;5HT2B::::8.8:C;ADA1A:::ant:8.72:DC;DRD2:::ant:8.55:DC;5HT7R:::ant:8.3:DC;HRH1:::ant:8.28:DC;DRD3:::ant:8.2:DC;ADA1B::RAT::8.1:C;DRD1:::ant:8.02:DC;H10::::7.82:C;HRH1::CAVPO::7.8:C;DRD4:::ant:7.49:DC;SC6A4::::7.28:C;5HT6R:::ant:7.21:DC;KCNH2::::6.92:C;HRH1::RAT::6.82:C;ADA2A:::ant:6.41:DC;5HT3A:::ant:6.4:DC;ADA2C::RAT::6.3:C;RORG::MOUSE::5.35:C;ACM1:::ant:5.29:DC;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ADA2C:::ant::D;ADA2B:::ant::D;ADA1B:::ant::D;5HT1E:::ant::D;5HT1D:::ant::D;5HT1B:::ant::D;DRD5:::ant::D|AOXA:::sub::D;CP3A4:::sub::D||
Methysergide|ok|5HT2B:::ant:9.45:DC;5HT2C:::ant:8.96:DC;5HT2B::RAT::8.84:C;5HT2A::RAT::8.84:C;5HT2A:::ant:8.8:DC;5HT7R::RAT::7.9:C;5HT7R:::ant:7.9:DC;5HT1A::RAT::7.51:C;5HT1B::RAT::7.5:C;DRD3::::7.23:C;5HT6R::::7.12:C;DRD2::::6.57:C;DRD1::::6.33:C;ADA2A::::6.21:C;SGMR1::::6.04:C;ADA2B::::5.66:C;AL1A1::::5.5:C;5HT1E:::bin::D;5HT1F:::bin::D;5HT1B:::bin::D;5HT1A:::ago::D|CP3A4:::sub::D||
Cabergoline|ok|5HT2B:::ago:8.85:DC;DRD1,DRD5:::ago::D;ADRB2:::bin::D;ADRB1:::bin::D;ADA1D:::bin::D;ADA1B:::bin::D;ADA1A:::bin::D;5HT7R:::ant::D;5HT2C:::ago::D;5HT1B:::ago::D;DRD1:::ago::D;DRD5:::ago::D;ADA2C:::ant::D;5HT1A:::ago::D;ADA2A:::ant::D;DRD4:::ago::D;5HT1D:::ago::D;ADA2B:::ant::D;5HT2A:::ago::D;DRD3:::ago::D;DRD2:::ago::D|CP3A4:::inh::D|MDR1:::sub::D|
Idoxuridine|ok_inv|KITH::::7.05:C;KITH::HHV1:::D;DNA|||
Dapsone|ok_inv|5HT6R::::6.74:C;LMNA::::5.85:C;DYR::PNECA::5.82:C;TSHR::::5.1:C;DHPS1::MYCLE:inh::D;DHPS2::MYCLE:inh::D|CP3A4:::sub:5.1:DC;CP2CI:::sub::D;PERM:::sub::D;CP2E1:::sub::D;CP3A7:::sub::D;CP2C9:::sub_ind::D;ARY2:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;PGH2:::sub::D;PGH1:::sub::D;FMO3:::sub::D;CP3A5:::sub::D||
Terconazole|ok|ADA2C::::7.21:C;SGMR1::::6.67:C;ADA2A::::6.43:C;ADA2B::::5.9:C;ACM1::::5.86:C;HS90A::::5.85:C;DRD3::::5.8:C;ACM4::::5.72:C;5HT2A::::5.63:C;LOX15::RABIT::5.61:C;5HT4R::CAVPO::5.61:C;CP51A::::5.52:C;ACM3::::5.51:C;ACM5::::5.5:C;5HT2C::::5.44:C;SC6A3::::5.36:C;ACM2::::5.34:C;ADA1A::RAT::5.27:C;SC6A4::::5.22:C;ADA1D::::5.15:C;AMPC::ECOLI::5.15:C;ADA1B::RAT::5.1:C;NR1I2::::5.05:C;NR1I2::RAT::5.04:C;CP51::CANAL:ant::D|||
Phenytoin|ok_vet|BLM::::8.66:C;ACM1::RAT::5.85:C;IMPA1::RAT::5.3:C;RORG::MOUSE::5.2:C;END4::ECOLI::5.1:C;GABAR;SCN8A:::inh::D;SCN2A:::inh::D;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1A:::inh::D;KCNH2:::inh::D;SCN3A;SCN1B;NR1I2;SCN1A:::inh::D;SCN5A:::inh::D|CP2C9:::duo:5.22:DC;CP2CI:::sub::D;NQO1:::sub::D;COMT:::sub::D;UD14:::sub::D;HYEP:::sub::D;CP2E1:::sub::D;CP2D6:::sub::D;CP2A6:::sub::D;CP1A2:::ind::D;UD19:::inh::D;UD16:::inh::D;UD11:::sub_ind::D;C11B1:::inh::D;CP3A7:::sub_ind::D;CP3A5:::sub_ind::D;CP3A4:::sub_ind::D;CP2B6:::sub_ind::D;CP2C8:::sub_ind::D;CP2CJ:::sub::D|MRP2:::sub::D;MDR1:::sub::D;SO1C1:::inh::D|THBG:::sub::D;ALBU
Medrysone|ok|GCR:::ago::D|CP3A5:::ind::D;CP3A4:::sub_ind::D||CBG
Doxycycline|ok_inv_vet|16S_ribosomal_RNA::Gut_flora:bin::D|CP3A4:::inh::D|ABCB5:::ind::D;S22A6:::inh::D|
Diethylstilbestrol|ok_inv|ESR2:::ago:10.7:DC;ESR1:::ago:10.22:DC;MK01::::6.5:C;AOXA::::6.34:C;ERR3:::ago:6.2:DC;SC6A3::::6.07:C;OPRD::::6.02:C;AA3R::::5.9:C;5HT2A::::5.86:C;AA1R::::5.78:C;OPRK::::5.74:C;5HT2B::::5.7:C;ADA2C::::5.66:C;OPRM::::5.63:C;LOX15::RABIT::5.53:C;DRD3::::5.52:C;NK2R::::5.5:C;SC6A2::::5.44:C;ACM1::::5.44:C;DRD1::::5.41:C;ACM3::::5.41:C;THAS::::5.36:C;DRD2::::5.35:C;GCR::::5.32:C;AA2AR::::5.3:C;ADA2A::::5.28:C;ADA2B::::5.27:C;ADA1D::::5.27:C;PGH1::::5.25:C;5HT6R::::5.22:C;SC6A4::::5.18:C;ADA1A::RAT::5.1:C;CLTR1::::5.05:C;KMT2A::::5.:C;SHBG;ANDR:::ant::D;NR1I2;NCOA2;ERR2;ERR1|CP3A4:::inh:5.:DC;CP2E1:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;CP19A:::inh::D;COMT:::sub::D|ABCG2:::inh:6.3:DC;ABCBB:::sub::D;SO2B1:::sub::D;SO1B1:::inh::D;MDR1:::sub::D|TTHY
Lymecycline|ok_inv|RS9::ECOLI:inh::D;RS4::ECOLI:inh::D|||
Clotrimazole|ok_vet|CP19A::::8.74:C;LMNA::::8.35:C;THAS::::7.85:C;CP2CJ::::7.8:C;KCNN4:::inh:7.15:DC;CP121::MYCTU::7.14:C;NR1I3::::7.1:C;CP17A::::7.09:C;CP51A::::6.89:C;CP51::MYCTU::6.7:C;CAC1C::::6.23:C;OPRM::::6.14:C;DRD3::::6.05:C;CP1A2::::5.9:C;GCR::::5.83:C;CCR4::::5.8:C;ACM4::::5.79:C;ACM1::::5.78:C;OPRD::::5.76:C;CXCR1::::5.7:C;ACM3::::5.68:C;MEN1::::5.65:C;V2R::::5.6:C;OPRK::::5.6:C;AA3R::::5.57:C;KCNH2::::5.52:C;SC6A4::::5.51:C;5HT2A::::5.5:C;NR1H4::::5.49:C;HRH1::::5.47:C;NK2R::::5.47:C;MDR1B::MOUSE::5.46:C;ADA2B::::5.43:C;DRD2::::5.39:C;ADA2A::::5.35:C;DRD1::::5.35:C;SC6A3::::5.35:C;ADRB2::::5.33:C;MDR1A::MOUSE::5.32:C;NPSR1::::5.3:C;HIF1A::::5.3:C;HRH2::::5.29:C;ACM2::::5.29:C;ADRB3::::5.27:C;I23O2::MOUSE::5.23:C;5HT6R::::5.23:C;KCNA3::::5.22:C;STRP::STRP1::5.21:C;P53::::5.2:C;RORG::MOUSE::5.2:C;ADRB1::::5.19:C;DRD4::::5.16:C;ACM1::RAT::5.15:C;AA2AR::::5.15:C;ADA1D::::5.13:C;5HT2B::::5.13:C;5HT2C::::5.12:C;AA1R::::5.11:C;ANDR::RAT::5.11:C;SC6A2::::5.1:C;AGAL::::5.1:C;NK1R::::5.06:C;FRIL::HORSE::5.05:C;5HT1A::RAT::5.:C;Ergosterol::CANAL:inh::D;HCAR2:::pag::D;NR1I2:::act::D;CP51::CANAL:ant::D|CP2C9:::inh:7.8:DC;CP3A4:::duo:7.8:DC;CP2C8:::inh:6.1:DC;CP2D6:::inh:6.05:DC;CP3A7:::ind::D;CP2E1:::inh::D;CP2A6:::inh::D;CP2B6:::duo::D|MDR1:::duo:5.89:DC;SO1B3:::ind::D;SO1B1:::inh::D;ABCBB:::inh::D|
Calcium_acetate|ok_inv|Phosphate:::bin::D|||
Sulfanilamide|ok|CAH13::MOUSE::7.49:C;CAH13::::7.49:C;CAH12::::7.43:C;CAH7::::7.15:C;CAH9::::6.62:C;CAH2::::6.62:C;CAN::CANAL::6.62:C;CAH::METTE::6.6:C;CAH1::::6.52:C;CYNT::HELPY::6.37:C;CAH2::BOVIN::6.07:C;CAH6::::6.03:C;CAH3::::6.01:C;TSHR::::6.:C;CAH4::BOVIN::5.52:C;CAH4::::5.52:C;CAH5B::::5.44:C;CAH14::::5.27:C;MTCA1::MYCTU::5.03:C;CAH15::MOUSE::5.02:C;DHPS::ECOLI:inh::D|CP3A4:::inh::D;CP2E1:::inh::D;CP2D6:::inh::D;CP2CJ:::inh::D||
Cycloserine|ok|HIF1A::::5.8:C;NMDZ1::RAT::5.64:C;TSHR::::5.4:C;MK01::::5.3:C;LMNA::::5.2:C;CP3A4::::5.:C;ALR::MYCAV:inh::D;DDLA::ECOLI:inh::D|DDC:::inh::D|S36A2|
Anagrelide|ok|PDE3A:::inh:7.3:DC;P2Y12::::5.98:C|CP1A2:::inh::D||
Carmustine|ok_inv|BLM::::7.85:C;AL1A1::::5.5:C;GSHR:::inh:5.09:DC;END4::ECOLI::5.:C;RNA;DNA|||
Sulfisoxazole|ok_vet|CP2CJ::::8.2:C;TSHR::::6.4:C;EDNRA::::6.11:C;EDNRA::RAT::6.11:C;MEN1::::5.15:C;DHPS::ECOLI:inh::D|CP2C9:::inh::D||
Metoprolol|ok_inv|ADRB1:::ant:7.8:DC;ADRB1::RAT::7.64:C;ADRB2::CAVPO::6.79:C;ADRB1:W134A:RAT::6.2:C;ADRB2:::ant:5.75:DC;ADRB1:S190A:RAT::5.6:C;ADRB1:Y356F:RAT::5.6:C;CP2J2::::5.31:C;ADRB1:Y356A:RAT::5.3:C;5HT1A::RAT::5.:C|CP3A4:::sub::D;CP2D6:::inh::D|MDR1:::sub::D;S22A2:::inh::D|ALBU:::bin::D
Crotamiton|ok||||
Dicoumarol|ok|NQO1:::inh:8.59:DC;GPR35::::7.41:C;LMNA::::7.3:C;PCSK7::::5.89:C;ALDR::RAT::5.39:C;MK01::::5.35:C;CP3A4::::5.3:C;AL1A1::::5.2:C;P53::::5.:C;CP2CJ::::5.:C;QOR:::inh::D;VKOR1:::inh::D|CP2C9:::sub:7.6:DC;CP2CB::RAT:inh::D;CP2C6::RAT:inh::D||ALBU
Cefmenoxime|ok|PBPA::CLOPE:inh::D;FTSI::ECOLI:inh::D|||
Ropinirole|ok_inv|DRD3:::ago:8.54:DC;DRD2:::ago:8.43:DC;DRD3::RAT::8.41:C;DRD4:::ago:8.11:DC;DRD2::RAT::7.12:C;5HT2A::::6.85:C;CP3A4::::6.5:C;5HT1A::::5.77:C;CP2D6::::5.5:C;DRD2::BOVIN::5.17:C;ADA1A,ADA1B,ADA1D,ADA2A,ADA2B,ADA2C:::ant::D|CP1A2:::sub::D||
Chlorotrianisene|inv_out|CP2CJ::::7.:C;LMNA::::6.55:C;TAU::::5.25:C;NPSR1::::5.1:C;HIF1A::::5.:C;ESR1:::ago::D|CP19A:::ind::D||
Isradipine|ok_inv|CAC1C:::inh:8.66:DC;CAC1C::RABIT::6.97:C;CAC1D::RAT::6.66:C;CP2C9::::5.44:C;CP2D6::::5.32:C;CP2C8::::5.3:C;CAC1S:::inh::D;CAC1D:::inh::D;CA2D2:::inh::D;CAC1H:::inh::D;CACB2:::inh::D;CA2D1:::inh::D|CP3A4:::inh:5.:DC|ABCBB:::sub::D|
Diatrizoate|ok_vet||||
Betazole|ok|LMNA::::5.95:C;HRH2:::ago::D|||
Topiramate|ok|CAH7::::9.06:C;CAH12::::8.42:C;CAH2:::inh:8.3:DC;CAN::CANAL::8.:C;CAH5A::::7.6:C;CAH5B::::7.6:C;CAH6::::7.35:C;CAH13::MOUSE::7.33:C;CAH13::::7.33:C;CAH4::BOVIN::7.27:C;CAH9::::7.24:C;CAH15::MOUSE::7.11:C;CAN::YEAST::6.96:C;CAH::METTE::6.92:C;CYNT::HELPY::6.76:C;CAH1:::inh:6.6:DC;MTCA2::MYCTU::6.32:C;MTCA1::MYCTU::6.21:C;CAH2::RAT::5.85:C;CAH14::::5.84:C;CAH4:::inh:5.31:DC;CAC1E:::ant::D;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4:::ant::D;CAH3:::inh::D;GRIK1,GRIK2,GRIK3,GRIK4,GRIK5:::ant::D;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A:::inh::D;GBRA1:::ago::D|CP3A4:::ind::D;CP2CJ:::inh::D|AAPK1,AAPK2,AAKB1,AAKB2,AAKG1,AAKG2,AAKG3:::ind::D;MDR1:::sub::D|ALBU:::bin::D
Cefmetazole|ok_inv|DACC::ECOLI:inh::D;DACA::ECOLI:inh::D;FTSI::ECOLI:inh::D;PBPB::ECOLI:inh::D;PBPA::ECOLI:inh::D;PBP2A::STAAU:inh::D||S15A2:::inh::D;S15A1:::inh::D|ALBU
Olmesartan|ok_inv|AGTR1::BOVIN::8.11:C;AGTR1:::ant::D||ABCBB:::sub::D;SO1B1:::sub::D;SO1B3:::sub::D;MRP2:::sub_ind::D|ALBU:::bin::D
Amsacrine|ok_inv|AOXA::RABIT::7.22:C;MTOR::::6.88:C;KCNH2:::inh:6.68:DC;TOP2A:::inh:6.14:DC;P53::::6.:C;TPO::::5.6:C;AOXA::RAT::5.52:C;AOXA::::5.49:C;HIF1A::::5.3:C;S22A1::::5.3:C;ACM1::RAT::5.2:C;CP2D6::::5.12:C;CP1A2::::5.1:C;ALBU;A1AG1;DNA:::itc::D||MDR1:::inh::D|
Theophylline|ok|AA1R:::ant:9.22:DC;AA2AR:::ant:9.22:DC;AA3R::::7.85:C;AA2BR::RAT::6.82:C;AA1R::RAT::6.15:C;LEF::BACAN::6.1:C;AA1R::BOVIN::5.61:C;AA2BR:::ant:5.57:DC;HIF1A::::5.5:C;AA2AR::RAT::5.17:C;AA1R::CAVPO::5.01:C;TTLL3;RIC3;PARP1;NOMO1;HM13;CPNE1;HDAC2:::act::D;PDE3A:::inh::D;PDE4A:::inh::D;PDE5A:::inh::D;PDE4B:::inh::D|CP2D6:::sub::D;CP1B1:::sub::D;CP1A1:::inh::D;CP2E1:::sub::D;ADA:::duo::D;CP1A2:::sub::D;CP3A4:::sub::D|S22A7:::inh::D|
Argatroban|ok_inv|THRB:::inh::D|CP3A5:::sub::D;CP3A4:::sub::D||A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Liothyronine|ok_vet|THA:::ago:10.24:DC;THB:::ago:10.1:DC;THB::RAT::8.74:C;AA1R::::6.62:C;NPSR1::::6.1:C;LMNA::::5.55:C;PCNA:::ant:5.44:DC;GBRP::RAT::5.15:C;MEN1::::5.1:C|UD11:::sub::D|LAT1;MDR1:::ind::D;MOT10:::inh::D;S22A8:::inh::D;SO4A1:::inh::D;SO1C1:::inh::D;NTCP:::sub::D;SO4C1:::sub::D;SO1B3:::sub::D;SO1B1:::sub::D;SO1A2:::sub::D|ALBU;THBG:::sub::D;TTHY
Disopyramide|ok|BLM::::6.25:C;THB::::5.5:C;A1AG2;KCNH2:::inh::D;KCND3:::inh::D;KCND2:::inh::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;SCN5A:::inh::D|CP1A2:::sub::D;CP3A4:::sub::D|S22A2:::inh:5.54:DC;S22A1:::inh::D|A1AG1
Lidocaine|ok_vet|AMPC::ECOLI::6.45:C;AL1A1::::6.05:C;SCN4A::::5.7:DC;A1AG2;A1AG1;EGFR:::ant::D;SCN5A:::inh::D;SCN9A:::inh::D;SCNAA:::inh::D|CP3A4:::sub:5.7:DC;CP2B6:::sub::D;CP2A6:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D;CP1A2:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP2D6:::inh::D|MDR1:::inh::D;S22A5:::inh::D|
Pamidronic_acid|ok|FPPS:::inh:7.25:DC;Hydroxylapatite:::ant::D|||
Clemastine|ok_inv|HRH1:::ant:10.31:DC;DRD3::::8.6:C;ACM4::::8.56:C;ACM5::::8.22:C;ACM3::::8.08:C;5HT2A::::8.04:C;ADA2C::::7.85:C;SGMR1::::7.85:C;ADA1D::::7.82:C;ADA1A::RAT::7.68:C;5HT2B::::7.64:C;5HT6R::::7.44:C;ADA1B::RAT::7.39:C;DRD2::::7.35:C;5HT2C::::7.28:C;ACM1::RAT::7.25:C;ADA2A::::7.16:C;ADA2B::::6.85:C;5HT1B::RAT::6.66:C;KCNH2::::6.49:C;HRH2::::6.44:C;SC6A3::::6.27:C;CP2CJ::::6.22:C;DRD1::::6.12:C;CP3A4::::5.6:C;SC6A2::::5.51:C;S22A1::::5.31:C;TPO::::5.:C|CP2D6:::inh:6.1:DC||
Acarbose|ok_inv|LYAG::RAT::6.8:C;SUIS::RAT::6.4:C;AMY1::::6.3:C;LYAG:::inh:5.35:DC;SUIS:::inh::D;AMYP:::inh::D;MGA:::inh::D|||
Venlafaxine|ok|LMNA::::8.7:C;SC6A4:::inh:8.42:DC;SC6A4::RAT::7.6:C;ADA1A::RAT::7.05:C;SC6A2:::inh:6.83:DC;SC6A3::RAT::6.44:C;SC6A3:::inh:5.44:DC|CP3A4:::sub::D;CP2D6:::inh::D|ABCG2:::ind::D;MDR1:::inh::D|
Conjugated_estrogens|ok|ESR1:::ago::D;ESR2:::ago::D|CP3A4:::sub::D;CP1A2:::inh::D;COMT:::sub::D|MRP3:::inh::D;MRP4:::inh::D;MRP1:::inh::D;SO1A2:::inh::D;NTCP:::inh::D;S22AA:::inh::D;S22A8:::inh::D;SO1C1:::inh::D;SO1B1:::inh::D;SO2B1:::sub::D;MDR1:::sub::D;S22A6:::sub::D;OSTA:::sub::D;OSTB:::sub::D;MRP2:::sub::D;SO4A1:::sub::D;ABCCB:::sub::D;SO1B3:::sub::D;S22AB:::sub::D;SO3A1:::sub::D;ABCG2:::sub::D|THBG:::ind::D;SHBG:::bin::D;ALBU:::bin::D
Travoprost|ok|PF2R:::ago::D|||
Amcinonide|ok|HIF1A::::8.89:C;NPSR1::::5.4:C;RORG::MOUSE::5.05:C;ANXA1:::ago::D;GCR:::ago::D|CP3A5:::ind::D;CP3A4:::sub_ind::D||
Atomoxetine|ok|SC6A2:::inh:8.69:DC;SC6A4:::bin:8.05:DC;SC6A4::RAT::7.37:C;SC6A3::RAT::6.15:C;SC6A3::::5.97:C;KCNH2::::5.68:C;OPRK:::pag::D;KCNJ3:::inh::D;NMDA:::inh::D|CP2D6:::sub:5.7:DC;CP2CJ:::sub::D||FCGR1:::bin::D;A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Bleomycin|ok_inv|DNLI3:::inh::D;DNA:::cli::D;DNLI1:::inh::D|BLMH:::sub::D||
Chlorambucil|ok|TSHR::::6.2:C;HIF1A::::5.3:C;LMNA::::5.15:C;NFKB1::::5.05:C;ALDR::RAT::5.03:C;TPO::::5.:C;DNA:::cov::D|GSTP1:::sub::D|SO1A2|
Etomidate|ok|GBRA1:::ago:5.92:DC;GBRB2::::5.46:C;GABAR:::aga::D;ADA2B:::ago::D|C11B2:::inh:10.:DC;C11B1:::inh:9.3:DC||GTR1:::inh::D
Raltitrexed|ok_inv|S19A1::::8.2:C;FOLR1::::7.82:C;FOLR2::::7.66:C;PCFT::::7.:C;TYSY:::inh:6.59:DC;TYSY::MOUSE::6.38:C;DRTS::TOXGO::6.32:C;TYSY::RAT::6.05:C;TYSY::ECOLI::5.64:C;TYSY::LACCA::5.1:C;FOLC:::ant::D|||
Etonogestrel|ok_inv|ESR1:::ago::D;PRGR:::ago::D|CP3A4:::sub::D||SHBG:::car:8.23:DC;ALBU:::car::D
Morphine|ok_inv|SGMR1::RAT::10.57:C;OPRM:::ago:9.85:DC;OPRM::RAT::9.85:C;OPRM::BOVIN::9.3:C;OPRM::CAVPO::9.06:C;OPRM::MOUSE::8.9:C;OPRK::CAVPO::8.74:C;OPRD::RAT::8.74:C;ADA2A::::8.52:C;OPRK:::ago:8.16:DC;OPRX::CAVPO::7.86:C;OPRD:::ago:7.81:DC;OPRK::RAT::7.57:C;OPRK::MOUSE::6.84:C;OPRD::MOUSE::6.81:C;LY96:::act::D|UD13:::sub::D;UD2B4:::sub::D;UDB15:::sub::D;UD18:::sub::D;UD11:::sub::D;UD2B7:::sub::D;CP3A4:::sub::D;CP2C8:::sub::D|MDR1:::sub::D|ALBU:::bin::D
Ropivacaine|ok|LMNA::::5.6:C;SCNAA:::inh::D|CP3A4:::sub::D;CP2B6:::sub::D;CP1A2:::sub::D||
Bupivacaine|ok_inv|SCN1A::::5.27:C;PE2R1;SCNAA:::inh::D|CP2D6:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D||
Dapiprazole|ok|ADA1D:::ant:8.39:DC;ADA1B::RAT::7.52:C;ADA1A::RAT::7.41:C;5HT2A::::6.76:C;5HT2C::::6.49:C;ADA2B::::6.28:C;5HT2B::::6.17:C;5HT1A::RAT::5.93:C;ADA1B:::ant::D;ADA1A:::ant::D|||
Penciclovir|ok|KITH::HHV1C:ind::D;DPOL::HHV11:inh::D|||
Tenofovir_disoproxil|ok_inv|DPOL::HBVD2:inh::D;Reverse_transcriptase_RNaseH::9HIV1:inh::D|KCRB,KCRM,KCRS,KCRU:::sub_ind::D;NDKA,NDKB:::sub::D;KAD4:::sub::D;KAD2:::sub::D|MDR1:::inh::D;MRP2:::sub::D;MRP4:::sub::D;MRP7:::sub::D;S22A8:::sub::D;S22A6:::sub::D|
Flucloxacillin|ok_inv|PBPA::CLOPE:inh::D|CP3A4:::sub_ind::D|ABCBB:::sub::D|
Tranexamic_acid|ok|PLMN:::inh:5.96:DC||S15A2|
Ertapenem|ok_inv|DACC::ECOLI:inh::D;PBPB::ECOLI:inh::D;PBPA::ECOLI:inh::D;DACB::ECOLI:inh::D;FTSI::ECOLI:inh::D;FTSI::HAEIN:inh::D;MRDA::ECOLI:inh::D;MRDA::HAEIN:inh::D|||
Desogestrel|ok|ESR1:::ago::D;PRGR:::ago::D|UD11:::ind::D;CP2C9:::sub::D;CP3A4:::sub::D||SHBG:::bin:6.6:DC;ALBU:::bin::D
Mitomycin|ok|DNA:::ant_cov::D|NCPR:::sub::D||
Talbutal|ok_ill|GABAR:::aga::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|||
Bexarotene|ok_inv|RXRA:::ago:8.57:DC;RXRB:::ago:8.23:DC;RARA::::8.22:C;RXRG:::ago:8.08:DC;RXRG::MOUSE::7.7:C;RXRB::MOUSE::7.68:C;RXRA::MOUSE::7.4:C;RXRA::RAT::7.4:C;RARB::::7.3:C;RARG::::6.89:C;CP26B::::5.23:C;MEN1::::5.:C|CP2C8:::inh::D;CP3A4:::sub_ind::D||
Ibutilide|ok|KCNH2:::inh:8.:DC;KCJ11:::inh::D;KCNH7:::inh::D;KCNH6:::inh::D;KCNK6:::inh::D;KCNK1:::inh::D;CCG1:::act::D;CA2D1:::act::D;CACB1:::act::D;CAC1C:::act::D|||
Vindesine|ok_inv|TBB1:::inh::D|CP3A4:::sub::D||
Chlorthalidone|ok|CAH7::::8.55:C;CAH12::::8.35:C;CAH5B::::8.05:C;CAH13::MOUSE::7.82:C;CAH9::::7.64:C;CAH2::::6.86:C;CAH4::::6.71:C;CAH1:::inh:6.46:DC;CAH5A::::6.04:C;CAH6::::5.87:C;CAH14::::5.38:C;TAU::::5.25:C;S12A1:::inh::D|||ALBU
Pentobarbital|ok_inv_vet|GBRP::RAT::5.77:C;NR1I2:::act::D;NMDA:::ant::D;GABAR:::aga::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2A6:::ind::D;CP2CJ:::sub::D;CP3A4:::ind::D||
Valproic_acid|ok_inv|PPARG;PPARD;PPARA;HDAC2:::inh::D;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A,SCN1B,SCN2B,SCN3B,SCN4B:::inh::D;SSDH:::inh::D;ODO1:::inh::D;HDAC9:::inh::D;ACDSB:::inh::D|UD11:::inh::D;UD19:::sub::D;UDB15:::sub::D;UD2B7:::sub::D;UD13:::sub::D;UD16:::sub::D;UD110:::sub::D;UD18:::sub::D;UD14:::sub::D;CP3A4:::inh::D;CP2CJ:::inh::D;CP1A2:::inh::D;PGH1:::sub::D;CP3A5:::sub::D;CP2C9:::inh::D;CP2B6:::sub::D;CP2A6:::sub_ind::D|SO2B1:::inh::D;S22A7:::sub::D;MOT1:::sub::D;S22A8:::inh::D;S22A5:::inh::D;S22A6:::inh::D|ALBU
Capreomycin|ok|TLYA::MYCTU:inh::D|||
Zolmitriptan|ok_inv|DRD2::RAT::10.4:C;DRD1::RAT::9.52:C;5HT1D:::ago:9.12:DC;5HT1B:::ago:8.82:DC;5HT1A:::ago:8.74:DC;ADA2C::RAT::8.15:C;5HT1F:::ago::D|AOFA:::sub::D;CP1A2:::sub::D||
Acetaminophen|ok|TSHR::::6.8:C;MYG::::5.64:C;CAH12::::5.39:C;CAH2::::5.21:C;CAH3::::5.15:C;CAH7::::5.04:C;CAH15::MOUSE::5.03:C;CAH1::::5.:C;TRPV1:::act::D;PGH1:::inh::D;PGH2:::inh::D;TEBP:::inh::D|GSTM1:::sub::D;GSTP1:::sub::D;FAAH1:::sub::D;ARY2:::inh::D;ST1A3:::sub::D;ST1A1:::sub::D;UDB15:::sub::D;UD19:::sub::D;UD11:::sub::D;UD16:::sub::D;CP2A6:::sub::D;CP2D6:::sub::D;CP3A4:::sub_ind::D;CP1A2:::sub::D;CP2E1:::sub::D|MDR1:::inh::D|ALBU:::bin::D
Gefitinib|ok_inv|EGFR:::ant:10.:DC;ERBB2:L858R:::9.7:C;EGFR:L858R::ant:9.03:DC;EGFR:G719S::ant:8.96:DC;EGFR:L861Q::ant:8.85:DC;EGFR:G719C::ant:8.7:DC;RIPK2::::8.42:C;ERBB2::::8.21:C;GAK::::8.15:C;EGFR:T790M::ant:7.4:DC;IRAK1::::7.16:C;HCK::::6.96:C;EGFR:L858R-T790M::ant:6.85:DC;ERBB4::::6.8:C;LYN::::6.8:C;ERBB2:T790M:::6.76:C;ABL1:Q252H:::6.64:C;M3K19::::6.62:C;FRK::::6.6:C;MKNK1::::6.54:C;HIPK4::::6.51:C;SIK2::::6.5:C;ABL1:Y253F:::6.44:C;MKNK2::::6.44:C;LCK::::6.4:C;ABL1:E255K:::6.4:C;SLK::::6.4:C;TBA1A::RAT::6.39:C;KC1E::::6.37:C;ABL1:H396P:::6.34:C;STK10::::6.33:C;ABL1::::6.32:C;MK14::::6.3:C;ABL1:M351T:::6.28:C;IRAK4::::6.27:C;SBK1::::6.25:C;EPHA6::::6.23:C;MP2K5::::6.22:C;CDK7::::6.21:C;CHK2::::6.2:C;ABL1:F317L:::6.11:C;MK10::::6.1:C;ERBB3::::6.1:C;PTK6::::6.01:C;BLK::::6.:C;M4K4::::6.:C;FLT3:D835Y:::6.:C;EPHB4::::6.:C;SRC::::5.96:C;FLT3:D835H:::5.96:C;KS6A4::::5.92:C;PIM3::::5.9:C;KPCD3::::5.9:C;CTRO::::5.89:C;EPHB1::::5.89:C;MK09::::5.85:C;ULK3::MOUSE::5.85:C;EPHA5::::5.82:C;IRAK3::::5.82:C;UFO::::5.8:C;MK06::::5.8:C;ABL2::::5.8:C;M4K5::::5.8:C;RET::::5.77:C;KIT:A829P:::5.74:C;MINK1::::5.74:C;EPHA8::::5.74:C;MYLK2::::5.72:C;VGFR2::::5.72:C;ST17A::::5.7:C;PIM1::::5.7:C;M3K3::::5.68:C;ACK1::::5.64:C;KPCD2::::5.6:C;KCC2D::::5.6:C;FGR::::5.59:C;PHKG2::::5.57:C;FLT3::::5.54:C;DCLK3::::5.54:C;FLT3:N841I:::5.52:C;MK04::::5.51:C;BRSK1::::5.5:C;KCC2G::::5.5:C;EPHB6::::5.49:C;KC1D::::5.49:C;M3K2::::5.48:C;MET:Y1235D:::5.46:C;KPCD1::::5.46:C;FLT3:R834Q:::5.46:C;PHKG1::::5.43:C;ST17B::::5.42:C;EPHA1::::5.4:C;LIMK1::::5.4:C;NLK::::5.38:C;KIT:D816V:::5.37:C;NUAK2::::5.34:C;ABL1:F317I:::5.33:C;FLT3:K663Q:::5.29:C;KIT:D816H:::5.26:C;EPHA3::::5.26:C;LTK::::5.26:C;DAPK3::::5.24:C;STK36::::5.24:C;TXK::::5.22:C;VGFR3::::5.2:C;DMPK::::5.16:C;TNIK::::5.16:C;PI42C::::5.12:C|CP2CJ:::inh::D;CP2C9:::inh::D;CP1A1:::inh::D;CP3A5:::sub::D;CP2D6:::inh::D;CP3A4:::inh::D|ABCG2:::inh:6.4:DC;MDR1:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Codeine|ok_ill|OPRM:::ago:6.98:DC;OPRM::MOUSE::5.:C;OPRD:::ago::D;OPRK:::ago::D|UD2B4:::sub::D;UD2B7:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D|S22A1:::inh::D|
Piperacillin|ok|PBP1B::STRR6:inh::D;PBP2A::STRR6:inh::D;PBP2::STRR6:inh::D;PBP3::STREE:inh::D||S22A8:::sub::D;S22A6:::inh::D|
Dihydroergotamine|ok_inv|5HT1A::RAT::9.42:C;5HT1B::RAT::9.42:C;ADA2A:::ago:9.41:DC;5HT6R::::8.83:C;ADA2C::::8.82:C;ADA2B::::8.75:C;DRD3::::8.74:C;ADA1A::RAT::8.69:C;5HT2A::::8.64:C;DRD2::::8.53:C;ADA2C::RAT::8.43:C;5HT2B:::ago:8.36:DC;ADA1B::RAT::8.35:C;ADA1D::::7.85:C;ADA1A::::7.55:C;5HT2C::::7.33:C;5HT4R::CAVPO::6.8:C;DRD1::::5.92:C;S47A1::::5.55:C;TAU::::5.5:C;5HT1B:::ago::D;5HT1D:::ago::D|CP3A4:::inh:5.52:DC|MDR1:::inh::D|
Amitriptyline|ok|ADA1A::RAT::10.7:C;HRH1::RAT::10.7:C;HRH1:::ant:9.26:DC;ACM4::::9.13:C;SC6A4:::inh:9.05:DC;ACM1,ACM2,ACM3,ACM4,ACM5:::lig:8.56,7.54,8.26,9.13,8.24:DC;ACM1::::8.56:C;5HT2C:::ant:8.5:DC;ADA2B::::8.43:C;5HT2A:::ant:8.36:DC;ACM3::::8.26:C;ACM5::::8.24:C;ADA2C::::8.07:C;SC6A2:::inh:7.66:DC;ACM2::::7.54:C;ADA1B::RAT::7.38:C;5HT3A::RAT::7.36:C;5HT2B::::7.35:C;ADA1D:::ant:7.28:DC;DRD3::::7.21:C;5HT6R:::ant:7.19:DC;DRD1::::7.05:C;ACM1::RAT::6.9:C;ADA2A:::duo:6.88:DC;DRD5::::6.77:C;DRD2::::6.71:C;SGMR1:::ago:6.36:DC;HRH2::CAVPO::6.18:C;HRH2:::inh:6.14:DC;RET::::6.:C;SCN9A::::6.:C;5HT1A::RAT::5.94:C;SCN5A::::5.8:C;5HT1B::RAT::5.77:C;SCN2A::::5.51:C;KCNH2,KCNH6,KCNH7:::inh:5.48,,:DC;KCNH2::::5.48:C;CAC1C::RAT::5.43:C;NFKB1::::5.3:C;SC6A3::::5.21:C;HCD2::::5.1:C;SC6A4::RAT::5.07:C;5HT2C::RAT:ant::D;KCNQ3:::inh::D;5HT1B:::bin::D;OPRM:::bin::D;5HT1D:::bin::D;5HT7R:::ant::D;ADA1B:::ant::D;HRH4:::bin::D;KCNA1:::inh::D;KCNQ2:::inh::D;ADA1A:::ant::D;NTRK2:::ago::D;NTRK1:::ago::D;OPRK:::ago::D;OPRD:::ago::D;5HT1A:::duo::D|CP2D6:::sub:5.1:DC;UD14:::sub::D;UDB10:::inh::D;CP2C8:::inh::D;CP2B6:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D;CP2CJ:::inh::D;CP1A2:::sub::D|MDR1:::sub::D|A1AG1:::bin::D;ALBU:::bin::D
Floxuridine|ok|TYSY::MOUSE::9.4:C;LMNA::::8.4:C;STRP::STRP1::6.16:C;TYSY|CP2C9:::inh::D;TYPH:::sub::D||THBG:::ind::D
Tolcapone|ok_out|COMT::RAT::8.66:C;COMT:::inh:6.9:DC;GPR35::::5.13:C|CP2C9:::inh::D||
Fluorometholone|ok_inv|GCR:::ago:8.8:DC;HIF1A::::8.:C;LYAG::::6.75:C;NR1I2::RAT::6.4:C;RORG::MOUSE::6.35:C;ANDR::RAT::6.07:C;NR1I2::::5.89:C;HD::::5.2:C|CP3A5:::ind::D;CP3A4:::sub_ind::D||CBG
Nitroprusside|ok_inv|ANPRA:::ago::D|CP1A1:::inh::D||
Calcium_glucoheptonate|ok||||
Hydromorphone|ok_ill|OPRM:::ago:9.55:DC;OPRK:::ago:8.55:DC;OPRD:::pag:7.42:DC|UD2B7:::sub::D;UD13:::sub::D;CP2C9:::sub::D||ALBU:::bin::D
Indomethacin|ok_inv|ANDR::::9.85:C;PGH1:::inh:8.7:DC;PGH1::MOUSE::8.7:C;PGH2::RAT::8.54:C;PGH1::SHEEP::8.4:C;PGH1::BOVIN::8.39:C;PGH2:::inh:8.23:DC;PGH1::RAT::8.22:C;PGH2::MOUSE::8.19:C;IL8::::7.3:C;PD2R2::::7.3:DC;AK1C3:::inh:7.:DC;THAS::::7.:C;PGH2::SHEEP::6.47:C;PTGDS::MOUSE::6.3:C;NPSR1::::5.8:C;ALDR::RAT::5.44:C;S22A6::RAT::5.38:C;NOS2::MOUSE::5.35:C;MTOR::::5.33:C;ALDR::BOVIN::5.3:C;ALDR::::5.22:C;HIF1A::::5.2:C;LOX5::::5.15:C;CP1A2::::5.:C;KDM4E::::5.:C;PPARA:::ago::D;LGUL:::inh::D;PPARG:::act::D;PTGR2:::inh::D;PA2GA:::inh::D|UD2B7:::inh::D;UD11:::inh::D;UD19:::sub::D;EST1:::sub::D;CP2C9:::sub::D;CP2CJ:::inh::D|S22A6:::inh:5.52:DC;S22A8:::inh:5.23:DC;ABCBB:::sub::D;SO1B1:::inh::D;S22A7:::sub::D;NTCP:::sub::D;S22AB:::inh::D;ABCCB:::inh::D;MRP2:::inh::D;SO1A2:::inh::D;MRP1:::inh::D;MDR1:::inh::D;MRP6:::inh::D;MRP4:::inh::D;MRP3:::inh::D|ALBU
Ethambutol|ok|EMBA::MYCTU:inh::D;EMBB::MYCTU:inh::D;EMBC::MYCTU:inh::D|||
Metformin|ok|LMNA::::8.46:C;GPDA:::inh::D;ETFD:::inh::D;AAKB1:::ago::D||S47A2:::sub::D;S29A4:::sub::D;S47A1:::sub::D;S22A3:::sub::D;S22A2:::inh::D;S22A1:::sub::D|
Ipratropium|ok_exp|ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D||S22A4:::sub::D;S22A5:::sub::D|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Methadone|ok|OPRM:::ago:8.39:DC;AOXA::RAT::7.52:C;OPRK::::6.29:C;OPRD:::ago:5.96:DC;KCNH2::::5.01:C;ACHB2:::ant::D;ACHA4:::ant::D;ACHA3:::ant::D;ACHA7:::ago::D;5HT3A:::ant::D;NMDA:::ant::D|CP2B6:::sub_ind:5.:DC;CP2C9:::sub::D;CP2CI:::sub::D;CP1A2:::sub::D;CP19A:::sub::D;CP2C8:::sub::D;CP2D6:::inh::D;CP3A7:::sub::D;CP2CJ:::sub::D;CP3A4:::duo::D|MDR1:::inh:5.12:DC|ALBU;A1AG1
Olanzapine|ok_inv|HRH1:::ant:10.06:DC;HRH1::RAT::9.52:C;5HT2A:::ant:8.84:DC;H10::::8.7:C;ACM1:::ant:8.68:DC;DRD2:::ant:8.68:DC;5HT2C:::ant:8.55:DC;5HT2A::RAT::8.4:C;DRD3::RAT::8.32:C;5HT6R:::ant:8.3:DC;5HT2B::::8.2:C;HRH1::CAVPO::8.2:C;DRD2::RAT::8.15:C;ADA1A:::ant:8.14:DC;DRD1,DRD5:::ant:8.,7.05:DC;ACM5::::8.:C;DRD1:::ant:8.:DC;5HT2B::RAT::7.92:C;ACM4:::ant:7.9:DC;ADA1B::RAT::7.84:C;DRD4:::ant:7.72:DC;DRD3:::ant:7.7:DC;DRD1::RAT::7.7:C;ACM1::RAT::7.66:C;ADA1A::RAT::7.6:C;ACM3:::ant:7.59:DC;ADA1D::::7.35:C;DRD4::RAT::7.3:C;ADA2C::::7.11:C;5HT7R::::7.1:C;DRD5:::ant:7.05:DC;ACM2:::ant:7.:DC;ADA2B::::7.:C;ADA2A::::6.85:C;KCNH2::::6.74:C;5HT3A:::ant:6.7:DC;ADA2C::RAT::6.5:C;ALR::::6.43:C;5HT1B::RAT::6.36:C;SC6A4::::6.26:C;5HT1A,5HT1B,5HT1D,5HT1E,5HT1F:::inh:6.21,6.,,,:DC;5HT1A::RAT::6.21:C;5HT1A::::6.21:C;ADA1B:::ant:6.:DC;5HT1B::::6.:C;LOX15::RABIT::5.56:C;MEN1::::5.35:C;LYAG::::5.25:C;MK01::::5.2:C;GBRA1,GBRA2,GBRA3,GBRA4,GBRA5,GBRA6,GBRG1,GBRG2,GBRG3:::inh::D;ADRB1,ADRB2,ADRB3:::inh::D|CP3A4,CP343,CP3A5,CP3A7:::inh::D;CP3A4:::inh::D;UD14:::sub::D;CP2C9:::inh::D;CP2CJ:::inh::D;FMO3:::sub::D;CP2D6:::inh::D;CP1A2:::sub::D|MDR1:::sub::D|A1AG1:::bin::D;ALBU:::bin::D
Atenolol|ok|AA3R::::8.75:C;LMNA::::8.3:C;ADRB1:::ant:6.82:DC;ADRB2::CAVPO::5.93:C;ADRB2:::ant:5.:DC;5HT1A::RAT::5.:C|CP2D6:::sub::D|ABCBB:::sub::D|ALBU:::sub::D
Nitrofural|ok_inv_vet|LMNA::::7.95:C;RORG::MOUSE::5.2:C;CITC::ECOLI:inh::D;MDH::ECOLI:inh::D;GSHR::ECOLI:inh::D;POXB::ECOLI:inh::D|XDH:::sub::D||
Pimecrolimus|ok_inv|MTOR:::pot::D;FKB1A:::pot::D|CP3A4:::inh::D||
Omeprazole|ok_inv_vet|ATP4A:::inh:6.6:DC;MCL1::::5.5:C;FAS::::5.47:C;ATP4B::PIG::5.42:C;RORG::MOUSE::5.35:C;KPYM::::5.15:C;PGDH::::5.:C;AHR:::ago::D|CP2CJ:::inh:5.6:DC;CP3A4:::duo:5.:DC;CP2D6:::inh::D;CP2CI:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP1B1:::ind::D;CP1A2:::duo::D;CP1A1:::sub_ind::D|MDR1:::inh::D;MRP3:::ind::D;ABCG2:::inh::D|
Pyrazinamide|ok_inv|TSHR::::7.7:C;Probable_fatty_acid_synthase_Fas_Fatty_acid_synthetase::MYCTU:inh::D|AOXA:::sub::D;XDH:::sub::D||
Metixene|ok|CHLE::HORSE::5.8:C;ACM3:::ant::D;ACM2:::ant::D;ACM5:::ant::D;ACM4:::ant::D;ACM1:::ant::D|||
Cetirizine|ok|HRH1:::ant:8.23:DC||MDR1:::inh::D|
Terfenadine|ok_out|HRH1:::ant:9.:DC;KCNH2:::inh:8.05:DC;5HT2B::::7.52:C;HRH1::CAVPO::7.45:C;5HT2A::::7.14:C;TAU::::6.95:C;CAC1C::RAT::6.85:C;SC6A3::::6.69:C;CAC1C::CAVPO::6.6:C;DRD3::::6.29:C;ADA2C::::6.26:C;5HT6R::::6.22:C;5HT2C::::6.19:C;CCR5::::6.07:C;NK2R::::6.05:C;CAC1C::::6.03:C;SCN5A::::6.01:C;LMNA::::6.:C;END4::ECOLI::5.9:C;MEN1::::5.9:C;DRD1::::5.87:C;ADA1B::RAT::5.73:C;SC6A2::::5.72:C;MDR1B::MOUSE::5.7:C;DRD2::::5.69:C;ADA1A::::5.63:C;TPO::::5.6:C;ACM1:::bin:5.54:DC;HD::::5.5:C;EGFR::::5.45:C;FYN::::5.21:C;RORG::MOUSE::5.2:C;MTOR::::5.13:C;ACM1::RAT::5.1:C;ACM2:::bin::D;ACM4:::bin::D;ACM5:::bin::D;ACM3:::ant::D|CP3A4:::duo:6.49:DC;CP2J2:::inh:5.95:DC;CP2C8:::inh::D;CP3A5:::sub::D;CP2D6:::inh::D;CP3A7:::sub::D|MDR1:::inh:5.96:DC;ABCBB:::sub::D|
Diltiazem|ok_inv|CAC1C::RAT::7.8:C;CAC1D::RAT::7.34:C;CAC1S::::6.42:C;CAC1C:::inh:6.35:DC;CAC1C::CAVPO::6.2:C;SCN1A::::5.05:C;CCG1:::inh::D|CP3A4:::inh:7.:DC;CP2C8:::sub::D;CP2D6:::sub::D;CP2CJ:::sub::D;CP3A7:::inh::D;CP3A5:::inh::D|MDR1:::inh::D|A1AG1:::bin::D;ALBU:::bin::D
Protriptyline|ok|AA3R::::8.96:C;SC6A2:::inh:8.85:DC;LMNA::::8.15:C;ACM1::RAT::6.8:C;CP3A4::::5.4:C;CP2D6::::5.4:C;NFKB1::::5.05:C;TPO::::5.:C;P53::::5.:C;SC6A4:::inh::D||MDR1:::inh::D|
Aminohippuric_acid|ok_inv|HIF1A::::5.3:C;AMPC::ECOLI::5.25:C;S22A6::MOUSE::5.03:C||S22A6:::inh:5.22:DC;S22A7:::sub::D;MOT1:::sub::D;SO1A2:::sub::D;MRP1:::sub::D;SO1B1:::inh::D;SO3A1:::inh::D;S22AB:::inh::D;S22A4:::inh::D;MRP2:::inh::D;S22A8:::inh::D;S22A5:::inh::D;S22A2:::inh::D|
Alfuzosin|ok_inv|ADA1B:::ant:8.55:DC;ADA1D:::ant:8.5:DC;ADA1D::RAT::8.46:C;ADA1B::RAT::8.31:C;ADA1A:::ant:8.09:DC;ADA1A::BOVIN::7.64:C;ADA1A::RAT::7.61:C;KCNH2:::inh::D|CP3A4:::sub::D||
Trimethadione|ok|CAC1G:::inh::D|CP2CJ:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP3A4:::sub::D;CP2E1:::sub::D||
Nitisinone|ok_inv|HPPD:::inh:7.43:DC;HPPD::PIG::7.4:C|||
Clobazam|ok_ill|GABAR:::aga::D|CP2D6:::inh::D;CP2CI:::sub::D;CP2B6:::sub::D;CP2CJ:::sub::D;CP3A4:::sub_ind::D|MDR1:::sub::D;S6A11;SC6A1|
Minoxidil|ok_inv|TSHR::::5.2:C;RENI;PGH1:::ind::D;KCNJ1:::ind::D|UD11:::sub::D||
Megestrol_acetate|ok_inv_vet|GCR:::ago:8.06:DC;ANDR::RAT::7.7:C;NPSR1::::5.5:C;HIF1A::::5.1:C;LMNA::::5.05:C;CP2C9::::5.:C;PRGR:::ago::D|CP3A4:::sub::D|MDR1:::inh::D|
Tioguanine|ok|PGH1::::6.22:C;HBB::::5.95:C;PAX8::::5.93:C;P53::::5.4:C;MK03::::5.26:C;DNA:::itc::D|HPRT:::sub::D|MRP4:::inh::D|
Methylergometrine|ok|5HT2A::::9.14:C;5HT2B::::9.1:DC;5HT6R::::8.93:C;5HT1A::RAT::8.63:C;5HT2C::::8.18:C;5HT1B::RAT::8.03:C;DRD3::::7.24:C;CP2D6::::6.7:C;ADA2B::::6.68:C;DRD2::::6.56:C;DRD1:::ant:6.27:DC;ADA2A::::6.22:C;AL1A1::::5.45:C;TAU::::5.3:C|CP3A4:::inh::D||
Buclizine|ok|HRH1:::ant::D;ACM1:::ant::D|||
Aztreonam|ok|PBPA::PSEAE::5.48:C;AMPC::CITFR:pot::D;PBPC::BACSU:inh::D|||
Chlorzoxazone|ok|LMNA::::7.4:C;TPO::::6.9:C;NOS1::RAT::5.55:C;TSHR::::5.1:C;NOS3::::5.06:C;KCMA1|CP1A2:::sub:6.4:DC;CP2D6:::sub::D;CP3A4:::inh::D;CP2A6:::sub::D;CP1A1:::sub::D;CP2E1:::inh::D||
Aminoglutethimide|ok_inv|CP19A:::inh:8.28:DC;CP19A::RAT::6.59:C;CP11A:::inh::D|CP2CJ:::ind::D;CP3A4:::ind::D||
Mefloquine|ok_inv|GLRA1::::5.6:C;KCNH2::::5.59:C;CP1A2::::5.2:C;LMNA::::5.05:C;P53::::5.:C;CP2D6::::5.:C;AA2AR:::ant::D;HBA:::ant::D;Fe_II_protoporphyrin_IX::PLAFA:ant::D|ACES:::inh::D;CP19A:::inh::D;CHLE:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Sulfadiazine|ok_inv_vet|LMNA::::6.75:C;Dihydropteroate_synthetase::PLAFA:inh::D|CP3A4:::sub::D;CP2C8:::sub::D;CP2C9:::inh::D||
Sapropterin|ok_inv|NOS1::::5.95:C;TPH1:::cof::D;TY3H:::cof::D;NOS3:::cof::D;PH4H:::cof::D|PGH2:::ind::D||
Vinorelbine|ok_inv|TBB5:::ant::D|CP3A4:::sub::D;CP2D6:::inh::D|MDR1:::sub::D|
Anidulafungin|ok_inv|FKS1::ASPNC:inh::D|||
Clozapine|ok|HRH1:::ant:9.4:DC;5HT2A::RAT::9.16:C;ACM1:::ant:9.01:DC;H10::::9.:C;ADA2C:::ant:8.94:DC;5HT2A:::ant:8.92:DC;ADA1B::RAT::8.85:C;5HT2B::RAT::8.74:C;ACM1::RAT::8.68:C;5HT2C:::ant:8.54:DC;HRH1::RAT::8.54:C;5HT2A::BOVIN::8.52:C;5HT2B::::8.5:C;BLM::::8.46:C;ADA1A:::ant:8.43:DC;HRH1::CAVPO::8.42:C;5HT6R:::ant:8.4:DC;5HT7R:::ant:8.26:DC;5HT7R::RAT::8.2:C;5HT1A:::ant:8.2:DC;ACM4:::ant:8.2:DC;DRD2:::ant:8.15:DC;DRD1:::ant:8.12:DC;5HT2C::RAT::8.1:C;DRD4::RAT::8.05:C;ACM5:::ant:8.02:DC;DRD4:::ant:8.:DC;ADA1B:::ant:8.:DC;ADA2B:::ant:7.96:DC;HRH4:::ant:7.92:DC;DRD2::RAT::7.82:C;ADA1A::RAT::7.82:C;ADA1D::::7.77:C;ACM3:::ant:7.77:DC;ADA2A::RAT::7.72:C;DRD3::RAT::7.65:C;ADA2A:::ant:7.62:DC;5HT2B::MOUSE::7.55:C;DRD5::RAT::7.52:C;5HT3A::MOUSE::7.49:C;5HT1A::RAT::7.41:C;ADA2C::RAT::7.4:C;DRD1::RAT::7.37:C;ACM2::RAT::7.34:C;5HT3A::RAT::7.28:C;DRD3:::ant:7.06:DC;ACM2:::ant:7.:DC;DRD2::BOVIN::6.85:C;AA3R::::6.81:C;ADA1A::BOVIN::6.8:C;DRD1::BOVIN::6.74:C;5HT3A:::ant:6.73:DC;KCNH2::::6.72:C;DRD5::::6.7:C;5HT1B::RAT::6.68:C;DRD2::CHLAE::6.6:C;SC6A4::::6.54:C;DRD2::MOUSE::6.54:C;DRD1::PIG::6.38:C;DRD3::CHLAE::6.33:C;HRH3::::6.2:C;NFKB1::::6.:C;5HT1B:::ant:6.:DC;5HT1E:::ant:6.:DC;5HT5A::::6.:C;LMNA::::5.95:C;SC6A2::::5.84:C;5HT1A::MOUSE::5.7:C;MEN1::::5.65:C;HRH2::::5.45:C;CAC1C::::5.44:C;IMPA1::RAT::5.35:C;AOXA::::5.29:C;SGMR1::::5.07:C;GSTP1;CALY;5HT1D:::ant::D|CP2D6:::inh:5.1:DC;CP1A1:::ind::D;UD14:::sub::D;FMO3:::sub::D;CP2C8:::sub::D;CP2A6:::sub::D;CP2CJ:::inh::D;CP3A4:::duo::D;CP2C9:::sub::D;CP1A2:::inh::D|MDR1:::sub::D|
Sucralfate|ok|PEPA5:::inh::D;FGF2:::ago::D;EGF:::ind::D;FIBA:::bin::D|||
Grepafloxacin|ok_out|PARC::HAEIN:inh::D;GYRA::HAEIN:inh::D|CP3A4:::sub::D;CP1A2:::inh::D|MRP2:::inh::D;S22A5:::inh::D;S22A2:::inh::D;S22A6:::sub::D;MRP1:::sub::D;MDR1:::inh::D|
Doxylamine|ok_vet|NR1I3;ACM1:::ant::D;HRH1:::ant::D|Q14097:::ind::D||
Levonorgestrel|ok_inv|PRGR:::mod::D;S5A1:::inh::D;ESR1;ANDR:::bin::D;SHBG:::inh::D;GCR:::bin::D|CP3A4:::sub::D;CP3A5:::sub::D||
Norepinephrine|ok|ADA1B::RAT::8.92:C;ADA2C::RAT::8.32:C;ADRB3:::ago:8.26:DC;ADA1A:::ago:8.04:DC;LMNA::::7.95:C;ADA1D::RAT::7.92:C;ADA2A:::ago:7.52:DC;ADRB1::RAT::7.28:C;ADA2B:::ago:7.21:DC;ADA2C:::ago:7.2:DC;ADA2B::RAT::7.11:C;ADRB2::CAVPO::6.67:C;ADA1B::MESAU::6.58:C;ADA1A::RAT::6.55:C;ADA1A::BOVIN::6.35:C;TYDP1::::6.3:C;ADA2C::MOUSE::6.19:C;APEX1::::6.1:C;TAU::::5.9:C;DRD2::::5.89:C;ADRB3::RAT::5.8:C;RECQ1::::5.65:C;ADRB1:::ago:5.59:DC;ADRB2:::ago:5.48:DC;BLM::::5.45:C;ADRB2::RAT::5.38:C;ADRB2::CANLF::5.3:C;ADA2A::MOUSE::5.24:C;ADRB2::BOVIN::5.22:C;VMAT1:::bin::D;VMAT2:::bin::D;PH4H:::inh::D;ADA1D:::ago::D;ADA1B:::ago::D||PO5F1:::sub::D;S22A1:::sub::D;S22A5:::inh::D;S22A3:::inh::D;S22A2:::inh::D;SC6A2:::sub::D|
Cidofovir|ok|DPOL::HCMVA:inh::D|TYPH:::inh::D|S22A6:::inh::D|
Mirtazapine|ok|HRH1:::ant:8.8:DC;5HT2A::RAT::8.7:C;5HT2C::RAT::8.26:C;ADA2C::::7.74:C;ADA2A:::ant:7.7:DC;5HT2C:::ant:7.41:DC;CP2CJ::::7.3:C;CP2C9::::7.3:C;5HT2A:::ant:7.16:DC;ADA2B::::6.65:C;5HT7R::::6.58:C;ADA1B::RAT::6.22:C;DRD2::RAT::5.84:C;5HT3A::::5.54:C;ADA1A,ADA1B,ADA1D:::ant:5.5,,:DC;ADA1A::::5.5:C;DRD1::RAT::5.38:C;5HT1A::::5.3:C;DRD3::::5.24:C;OPRK:::ago::D;5HT3_serotonin_receptor:::ant::D|CP2D6:::sub:6.3:DC;CP1A2:::sub::D;CP3A4:::inh::D|SC6A4:::inh::D|
Meprobamate|ok_ill|LMNA::::6.35:C;GABAR:::aga::D;GBRA6:::ago::D;GBRA5:::ago::D;GBRA4:::ago::D;GBRA3:::ago::D;GBRA2:::ago::D;GBRA1:::ago::D|||
Thiethylperazine|ok_out|PDR5::YEAST::5.64:C;DRD4:::ant::D;DRD1:::ant::D;DRD2:::ant::D|||
Timolol|ok|ADRB2::CAVPO::9.78:C;ADRB2:::ant:9.7:DC;ADRB1:::ant:8.82:DC;ADRB1::RAT::8.5:C;ADRB1:W134A:RAT::8.1:C;ADRB1:Y356F:RAT::7.8:C;ADRB1:S190A:RAT::7.5:C;ADRB3::::6.47:C;5HT1A::RAT::6.21:C;ADRB1:Y356A:RAT::6.2:C;ACM1::RAT::5.3:C;NFKB1::::5.:C;ENLYS::BPT4:::D|CP2D6:::sub:5.1:DC;CP2CJ:::sub::D|MDR1:::sub::D|
Treprostinil|ok_inv|PI2R:::ago::D;PPARD:::ago::D;P2Y12:::ago::D|CP2C9:::sub::D||
Colestipol|ok|Bile_acids:::bin::D|||
Trihexyphenidyl|ok|ACM4:::ant:9.12:DC;ACM1:::ant:8.87:DC;ACM3:::ant:8.5:DC;ACM5:::ant:8.06:DC;ACM2:::ant:7.92:DC;SGMR1::::7.35:C;CP2D6::::5.61:C|||
Palonosetron|ok_inv|5HT3A:::ant:10.5:DC;KCNH2::::5.7:C|CP1A2:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D||
Dydrogesterone|ok_out|PRGR:::ago::D|CP3A4:::sub::D||
Mexiletine|ok_inv|5HT2B::::6.14:C;SCN2A::::5.54:C;KCNH2::::5.:C;AHR:::ago::D;SCN5A:::inh::D|CP3A4:::sub::D;CP2E1:::sub::D;CP2B6:::sub::D;CP2D6:::sub::D;CP1A2:::inh::D||
Dexrazoxane|ok_out|TOP2B;TOP2A:::inh::D|||
Amlodipine|ok|CAC1C::RAT::8.7:C;ADA2A::::6.65:C;ADA2C::::6.58:C;KCNK2::::6.4:C;CAC1C::CAVPO::6.24:C;CAC1C:::inh:5.92:DC;5HT6R::::5.87:C;ADA1A::::5.63:C;SC6A3::::5.36:C;ADA1D::::5.27:C;ADA1B::::5.1:C;A0A024R8I1,CAC1B::,HUMAN:inh::D;CAC1I:::inh::D;ASM:::inh::D;CAH1:::inh::D;CA2D3:::inh::D;CACB1:::inh::D;CAC1B:::inh::D|CP2D6:::inh::D;CP2C8:::inh::D;CP3A5:::inh::D;CP2B6:::inh::D;CP1A1:::inh::D;CP3A4:::sub::D|MDR1:::inh::D|
Tacrine|ok_out|CHLE:::inh:10.57:DC;CLAT::RAT::9.82:C;CHLE::HORSE::8.92:C;ACES::ELEEL::8.7:C;ACES:::inh:8.5:DC;ACES::TETCF::8.09:C;A4::::7.91:C;ACES::MOUSE::7.74:C;ACES::BOVIN::7.57:C;AOFA::RAT::7.4:C;ACHE::::7.36:C;ACES::RAT::7.34:C;HNMT::RAT::6.96:C;ACM2::MOUSE::6.66:C;CP2D6::::6.52:C;SC6A2::::6.29:C;S22A2::::6.17:C;S47A1::::5.96:C;ADA1A::RAT::5.95:C;ACM1::MOUSE::5.7:C;ACM2::RAT::5.68:C;NMDZ1::::5.31:C;ACM2::::5.24:C;ACM1::RAT::5.23:C;ACM2::PIG::5.2:C;SC6A4::RAT::5.12:C;EST1|CP1A2:::sub:6.3:DC|MDR1:::sub::D|
Oxyphencyclimine|ok|ACM3:::ant::D;ACM1:::ant::D;ACM2:::ant::D|||
Triamterene|ok|ACM1::RAT::8.66:C;LMNA::::7.35:C;TSHR::::6.9:C;NFKB1::::6.65:C;PGDH::::6.15:C;KDM4E::::5.95:C;HCD2::::5.9:C;AL1A1::::5.5:C;PTR1::LEIMA::5.47:C;CASP1::::5.44:C;CYSP::TRYCR::5.4:C;JAK2::::5.34:C;LEF::BACAN::5.3:C;END4::ECOLI::5.25:C;SMN::::5.2:C;CATG::::5.13:C;LOX12::::5.05:C;HIF1A::::5.:C;CASP7::::5.:C;RORG::MOUSE::5.:C;CP2D6::::5.:C;AGAL::::5.:C;SCNND:::inh::D;SCNNB:::inh::D;SCNNA:::inh::D;SCNNG:::inh::D|CP1A2:::sub:5.3:DC||
Valrubicin|ok|TOP2A:::inh::D;DNA:::itc::D|||
Procyclidine|ok|NMDZ1::::5.77:C;HRH1::RAT::5.17:C;ACM3:::ant::D;ACM4:::ant::D;ACM2:::ant::D;ACM1:::ant::D|||
Phenylephrine|ok|ADA1B:::ago:9.07:DC;ADA1A::BOVIN::8.05:C;ADA1A:::ago:7.26:DC;ADA2C::RAT::7.11:C;ADA1D::RAT::6.81:C;HIF1A::::6.6:C;ADA2A::::6.51:C;ADA2C::::6.47:C;ADA1A::RAT::6.01:C;ADA1B::MESAU::5.9:C;ADA1B::RAT::5.7:C;NFKB1::::5.45:C;ADRB1::::5.22:C;ADA1D:::ago::D|CP1A2:::ind::D;ST1A3:::sub::D;AOFB:::sub::D;AOFA:::sub::D||
Carbimazole|ok_inv|LMNA::::5.05:C;PERT:::inh::D|CP19A:::inh::D||
Digoxin|ok|LEF::BACAN::7.5:C;SO1A4::RAT::7.43:C;RORG::::6.96:C;P53::::6.8:C;AT1A2::RAT::6.66:C;AT1A1:::inh:6.54:DC;PAX8::::6.38:C;AT1A1::CANLF::6.3:C;LMNA::::6.25:C;RORG::MOUSE::5.85:C;STAT3::::5.73:C;RECQ1::::5.4:C|CP11A:::inh::D|SO1B1:::inh:5.49:DC;OSTB:::sub::D;OSTA:::sub::D;SO1A2:::sub::D;ABCBB:::sub::D;SO4C1:::sub::D;MDR1:::duo::D|
Sulpiride|ok_inv|CAH6::::9.1:C;DRD2::RAT::8.82:C;BLM::::8.8:C;CAH7::::8.44:C;CAH12::::8.41:C;DRD2:::ant:8.12:DC;DRD3:::ant:8.1:DC;CAH5B::::7.74:C;CAH9::::7.51:C;CAH2:::inh:7.4:DC;CAN::CANAL::7.4:C;CAH15::MOUSE::7.14:C;CAN::YEAST::6.91:C;CAH5A::::6.76:C;CYNT::HELPY::6.75:C;DRD2::CANLF::6.7:C;MTCA2::MYCTU::6.58:C;CAH4::BOVIN::6.21:C;ADA2A::::6.12:C;CAH1::::5.92:C;DRD5::RAT::5.8:C;DRD4::::5.68:C;MTCA1::MYCTU::5.64:C;TAU::::5.05:C;CAH3:::inh::D|CHLE:::inh::D||
Profenamine|ok|ACES::::6.59:C;CHLE::HORSE::6.14:C;ACM2:::ant::D;NMD3A:::ant::D;ACM1:::ant::D|CHLE:::inh:7.7:DC||
Nimodipine|ok_inv|LMNA::::8.74:C;CAC1C:::inh:6.96:DC;CAC1C::CAVPO::6.52:C;NR1I2::::6.41:C;TRPA1::MOUSE::6.1:C;CP2C9::::6.:C;CNR1::::5.86:C;NPSR1::::5.8:C;CP2CJ::::5.66:C;CP2J2::::5.47:C;CP1A2::::5.14:C;AA3R::::5.07:C;NR1H4::::5.05:C;AHR:::ago::D;MCR:::ant::D;CACB4:::inh::D;CACB3:::inh::D;CACB2:::inh::D;CACB1:::inh::D;CAC1S:::inh::D;CAC1F:::inh::D;CAC1D:::inh::D|CP3A4:::sub:5.75:DC||
Beclomethasone_dipropionate|ok_inv|AMPC::ECOLI::5.25:C;GCR:::ago::D|CP3A4:::sub_ind::D;CP3A5:::ind::D|SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::sub_ind::D|CBG:::bin::D
Carisoprodol|ok|LMNA::::8.25:C;ACM1::RAT::7.:C;TSHR::::6.2:C;TYDP1::::6.1:C;GBRA3:::mod::D;GBRA5:::mod::D;GBRG2;GBRB2:::mod::D;GBRA1:::ago::D|CP2CJ:::sub::D||
Progesterone|ok_vet|PRGR:::ago:10.:DC;MCR:::duo:9.41:DC;ESR1::RAT::8.41:C;PRGR::RABIT::8.22:C;ANDR:::ago:8.07:DC;FABPL::RAT::7.57:C;GCR:::pag:7.52:DC;ANDR::MOUSE::7.43:C;CBG::::7.38:C;SHBG:::bin:6.94:DC;ANDR::RAT::6.84:C;SGMR1::RAT::6.62:C;SGMR1::::6.59:C;SGMR1::CAVPO::6.18:C;S22A2::RAT::5.8:C;S5A1::RAT::5.8:C;GPBAR::::5.56:C;ERG2::YEAST::5.35:C;ACM1::RAT::5.25:C;LMNA::::5.2:C;TSHR::::5.:C;TPO::::5.:C;NPSR1::::5.:C;ESR2:::duo::D;A1AG1:::bin::D;OPRK:::ago::D;ESR1:::duo::D|CP3A4:::sub_ind:5.4:DC;CP2C9:::inh:5.26:DC;CP2D6:::sub::D;CP2A6:::ind::D;CP1B1:::sub::D;CP1A1:::sub::D;CP2CJ:::inh::D;CP3A7:::inh::D;CP3A5:::sub::D;CP17A:::inh::DC|S22A1:::inh:5.52:DC;S22A3:::inh:5.37:DC;SO1B3:::ind::D;ABCG2:::duo::D;SO1B1:::inh::D;NTCP:::inh::D;MRP1:::inh::D;ABCBB:::inh::D;S22A2:::inh::D;MDR1:::duo::D|
Phenylpropanolamine|ok_vet_out|ADA2A,ADA2B,ADA2C;ADRB2:::ago::D;ADRB1:::ago::D;DRD1:::pag::D|AOFA:::inh::D||
Sorafenib|ok_inv|VGFR2:::ant:10.68:DC;RAF1:::inh:9.:DC;DDR1::::8.82:C;FLT3:::ant:8.7:DC;HIPK4::::8.57:C;EGFR::::8.53:C;BRAF:::inh:8.52:DC;VGFR3:::ant:8.52:DC;PGFRB:::ant:8.4:DC;FLT3:K663Q::ant:8.35:DC;FGFR1:::inh:8.33:DC;RET:::inh:8.22:DC;M3K20::::8.2:C;DDR2::::8.18:C;RET:M918T::inh:8.13:DC;KIT:::ant:8.:DC;FLT3:N841I::ant:7.96:DC;HYES::::7.92:C;KIT:V559D::ant:7.8:DC;MK14::::7.8:C;FLT3:R834Q::ant:7.77:DC;KIT:V559D-T670I::ant:7.74:DC;VGFR1:::inh:7.74:DC;MK03::::7.74:C;CSF1R::::7.72:C;KIT:A829P::ant:7.7:DC;RET:V804M::inh:7.66:DC;KIT:L576P::ant:7.6:DC;BRAF:K97R::inh:7.58:DC;FLT3:D835H::ant:7.52:DC;BRAF:V600E::inh:7.42:DC;RET:V804L::inh:7.41:DC;MK15::::7.34:C;5HT2B::::7.25:C;LCK::::7.22:C;PGFRA::::7.21:C;TIE1::::7.17:C;ABL1::::7.1:C;CDK8::::7.1:C;FLT3:D835Y::ant:7.09:DC;M3K19::::7.:C;MK01::::6.96:C;CDKL2::::6.89:C;MKNK2::::6.89:C;MUSK::::6.89:C;ABL1:Q252H:::6.89:C;CDK7::::6.85:C;STK10::::6.85:C;UFO::::6.8:C;ABL1:T315I:::6.8:C;MP2K5::::6.72:C;AURKB::::6.7:C;MK11::::6.7:C;AURKC::::6.68:C;CDPK1::PLAF7::6.66:C;ABL1::MOUSE::6.65:C;MKNK1::::6.64:C;ABL1:M351T:::6.64:C;EPHB6::::6.62:C;KIT:V559D-V654A::ant:6.62:DC;EPHA6::::6.62:C;CDK19::::6.6:C;KC1A::::6.6:C;TNI3K::::6.55:C;KIT:D816V::ant:6.51:DC;M4K5::::6.5:C;EPHA5::::6.44:C;HIPK3::::6.41:C;SRC::::6.41:C;NTRK3::::6.4:C;PLK4::::6.4:C;KS6B1::::6.4:C;LYN::::6.4:C;TAOK1::::6.4:C;ABL1:Y253F:::6.38:C;5HT2C::::6.38:C;KIT:D816H::ant:6.37:DC;FRK::::6.36:C;CDKL3::::6.31:C;HIPK2::::6.3:C;ABL1:H396P:::6.28:C;HCK::::6.28:C;TAOK2::::6.27:C;LIMK1::::6.2:C;NTRK2::::6.2:C;NLK::::6.19:C;EPHA7::::6.17:C;M3K7::::6.16:C;ABL1:F317L:::6.11:C;EPHA2::::6.1:C;AURKA::::6.1:C;BLK::::6.1:C;EPHA8::::6.02:C;SLK::::6.:C;HIPK1::::5.96:C;5HT1A::::5.93:C;FGFR3::::5.9:C;RIPK2::::5.89:C;MYLK2::::5.89:C;ABL2::::5.89:C;EPHA4::::5.89:C;CDK17::::5.8:C;MINK1::::5.8:C;NTRK1::::5.8:C;EPHB1::::5.77:C;ABL1:F317I:::5.77:C;EPHB4::::5.74:C;EPHA3::::5.72:C;EPHB2::::5.72:C;5HT2A::::5.71:C;DYRK3::::5.7:C;TIE2::::5.68:C;TNK1::::5.64:C;STK33::::5.62:C;VGFR2::DANRE::5.59:C;FGFR2::::5.57:C;TAOK3::::5.57:C;CDK15::::5.54:C;CDK14::::5.54:C;CSK::::5.54:C;EPHA1::::5.51:C;MEN1::::5.5:C;5HT5A::::5.48:C;ABL1:E255K:::5.47:C;TTK::::5.46:C;MERTK::::5.44:C;MK09::::5.44:C;STK36::::5.42:C;CDK3::::5.42:C;KCC2B::::5.4:C;M4K4::::5.32:C;M4K1::::5.32:C;SRPK1::::5.3:C;INSR::::5.28:C;FGFR3:G697C:::5.23:C;CTRO::::5.21:C;CDK5::::5.21:C;5HT6R::::5.21:C;MK13::::5.18:C;TGFR2::::5.16:C;MYO3B::::5.15:C;5HT7R::::5.15:C;JAK3::::5.14:C;KS6A6::::5.12:C;CLK1::::5.12:C;MK12::::5.12:C;FGR::::5.11:C;TNIK::::5.1:C;IRAK1::::5.1:C;FYN::::5.08:C;CDK2::::5.06:C;RORG::MOUSE::5.05:C;LIMK2::::5.02:C;MYLK3::::5.02:C;SRMS::::5.01:C|UD11:::inh::D;UD19:::inh::D;CP2D6:::inh::D;CP2CJ:::inh::D;CP1A2:::sub::D;CP2C8:::inh::D;CP2B6:::inh::D;CP3A4:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP2C9:::inh::D|SO1B1:::inh::D;RBP1:::sub::D;MDR1:::inh::D;MRP2:::inh::D;MRP4:::inh::D;ABCG2:::inh::D|
Zoledronic_acid|ok|FPPS:::inh:10.15:DC;CAH2::::7.21:C;CAH14::::7.04:C;GGPPS::YEAST::6.59:C;CAH12::::6.5:C;LMNA::::6.2:C;ISPA::ECOLI::5.96:C;GGPPS:::inh:5.57:DC;CAH9::::5.27:C;MMP2::::5.15:C;Hydroxylapatite:::ant::D||MRP1:::sub::D|
Griseofulvin|ok_inv_vet|TSHR::::5.1:C;K1C12;TBA::CANAX:inh::D;TBB::CANAX:inh::D|CP3A4:::ind::D;CP1A2:::ind::D||
Nisoldipine|ok|CAC1C:::inh:8.52:DC;CAC1C::CAVPO::7.1:C;CP1A2::::6.:C;AA2AR::::5.64:C;AA3R::::5.4:C;NR1I2::::5.1:C;LMNA::::5.1:C;CAC1S:::inh::D;CAC1D:::inh::D;CACB2:::inh::D;CA2D1:::inh::D|CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|
Eszopiclone|ok_inv|GBRA1:::pot:7.3:DC;GBRA4::::6.99:C;GBRB2::::6.94:C;GBRA5:::ago::D;GBRA3:::ago::D;GABAR:::aga::D;GBRA2:::ago::D|CP2C8:::sub::D;CP3A4:::sub::D||
Ceruletide|ok|CCKAR:::ind::D|||
Alprazolam|ok_ill_inv|GBRP::RAT::8.48:C;GBRA5:::lig:8.:DC;GBRA2:::lig:7.92:DC;LMNA::::7.9:C;GBRA1:::lig:7.43:DC;GBRA3:::lig:7.16:DC;RORG::MOUSE::5.7:C;BRD4::::5.61:C;GBRA4:::lig::D;GABAR:::aga::D;TSPO:::lig::D;GBRA6:::lig::D|CP2C9:::sub::D;CP3A5:::sub::D;CP3A7:::sub::D;CP3A4:::sub::D||A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Dexbrompheniramine|ok|HRH1:::ant::D|||
Gentian_violet_cation|ok|DNAS1::::6.46:C;DNA:::itc::D||S22A1|
Ardeparin|ok_out|ANT3:::pot::D;HEP2:::ago::D|||
Loxapine|ok|5HT2A:::ant:8.62:DC;DRD4:::bin:8.31:DC;5HT2A::RAT::8.22:C;5HT6R:::bin:7.82:DC;ADA1B::RAT::7.74:C;DRD2::RAT::7.68:C;DRD2:::ant:7.68:DC;DRD3:::bin:7.66:DC;5HT7R::RAT::7.37:C;HRH4:::bin:6.66:DC;5HT2C::RAT::6.:C;HRH1::RAT::6.:C;ACM1:::bin:5.26:DC;SC6A3:::bin::D;SC6A2:::bin::D;SC6A4:::bin::D;HRH2:::bin::D;HRH1:::bin::D;DRD5:::bin::D;DRD1,DRD5:::bin::D;ACM5:::bin::D;ACM4:::bin::D;ACM3:::bin::D;ACM2:::bin::D;ADRB1:::bin::D;ADA2C:::bin::D;ADA2B:::bin::D;ADA2A:::bin::D;ADA1B:::bin::D;ADA1A:::bin::D;5HT7R:::bin::D;5HT5A:::bin::D;5HT3A:::bin::D;5HT1E:::bin::D;5HT1D:::bin::D;5HT1B:::bin::D;5HT1A:::bin::D;5HT2C:::ant::D;DRD1:::ant::D|||
Remoxipride|ok_out|DRD2:::ant:8.92:DC;SGMR1:::ant:7.26:DC;DRD2::CHLAE::6.06:C;DRD2::RAT::5.85:C;DRD5::RAT::5.8:C;HIF1A::::5.7:C;DRD4:::ant:5.41:DC;5HT1A::::5.4:C;DRD3::CHLAE::5.34:C;5HT2A;DRD3:::ant::D|CP2D6:::sub:6.7:DC||
Mupirocin|ok_inv_vet|SYIC::::9.1:C;SYI::THET8::6.6:C;STRP::STRP1::6.37:C;SYI1::STAAU:inh::D|||
Carbamoylcholine|ok|ACM4::::9.4:DC;ACM1::RAT::8.89:C;ACM2:::ago:8.42:DC;ACM2::RAT::8.4:C;ACM2::MOUSE::8.1:C;ACES::MOUSE::8.1:C;ACM1::MOUSE::7.7:C;ACM3::::7.15:DC;ACM1:::ago:6.77:DC;ACHA2::RAT::6.68:C;ACM4::RAT::6.64:C;ACM5::::6.44:C;ACHA3::RAT::6.35:C;ACM3::RAT::6.32:C;ACHA4::RAT::6.23:C;AMPC::ECOLI::5.3:C;ACHA::TETCF::5.12:C;ACM3::MOUSE::5.:C;ACES;ACHA2:::ago::D|PA24A:::ind::D||
Rosiglitazone|ok_inv|AGTRA::RAT::9.64:C;PPARG:::ago:9.:DC;LMNA::::8.66:C;PPARA::::8.4:DC;PPARG::MOUSE::7.52:C;CISD1::::7.51:C;AOFB::::6.08:C;CISD1::RAT::5.96:C;THAS::::5.45:C;PPARD::::5.44:DC;CAH2::::5.39:C;AOFB::RAT::5.24:C;RXRG;RXRB;RXRA;ACSL4:::inh::D|CP3A4:::sub:5.1:DC;CP2D6:::inh::D;CP2A6:::inh::D;CP1A2:::inh::D;PGH1:::sub::D;CP2C9:::sub::D;CP2C8:::inh::D|ABCBB:::sub:5.19:DC;SO1B1:::inh::D|ALBU:::sub::D
Pramipexole|ok_inv|DRD3::RAT::9.68:C;DRD4:::ago:9.31:DC;DRD3:::ago:9.14:DC;DRD2::BOVIN::8.8:C;DRD2::RAT::8.77:C;DRD2:::ago:8.3:DC;5HT2A::::5.93:C;ADA2A:::ago::D;5HT1A:::ago::D||S22A3;S22A1:::sub::D;S22A2:::sub::D|
Acetohexamide|ok_out|THB::::8.6:C;BLM::::8.55:C;TSHR::::8.2:C;KCNJ1:::inh::D|CP2C9:::sub::D;CBR1:::sub::D||ALBU
Ampicillin|ok_vet|AMPC::ECOLI::6.25:C;TIE2;PBP2::STRR6:inh::D;PBPA::STRR6:inh::D;PBP3::STREE:inh::D;PBP1B::STRR6:inh::D;PBP2A::STRR6:inh::D||MOT1;S22A5:::inh::D;S15A2:::inh::DC;S15A1:::inh::DC|ALBU
Metocurine_iodide|ok_out|ACHA2:::ant::D|||
Phenoxymethylpenicillin|ok_vet|S15A1;PAC::LYSSH:::D;DACB::ECOLI:::D;MecA::STAAU:inh::D;PBPA::CLOPE:::D|||
Secobarbital|ok_vet|MMP9::::5.58:C;NMDA:::ant::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2CJ:::ind::D;CP1A2:::ind::D;CP2C8:::ind::D;CP2C9:::ind::D||
Miglustat|ok|LYAG::::7.:C;GBA2::MOUSE::6.85:C;GBA2::::6.64:C;SUIS::::6.3:C;SUIS::RAT::6.24:C;LYAG::RAT::5.68:C;MGA::::5.68:C;LYAG::MOUSE::5.05:C;GDE::::5.:C;CEGT:::inh::D|||
Promazine|ok_vet|HRH1:::ant:9.4:DC;ADA1A::RAT::8.43:C;ADA1B::RAT::8.34:C;ADA1D:::ant:8.21:DC;5HT2A:::ant:8.17:DC;ADA2B::::8.07:C;SC6A2::::7.89:C;ADA2C::::7.43:C;TSHR::::7.4:C;ACM4:::ant:7.38:DC;ACM5:::ant:7.34:DC;SC6A4::::7.34:C;5HT2C:::ant:7.28:DC;DRD3::::7.16:C;ACM3:::ant:7.06:DC;SGMR1::::6.94:C;ACM1:::ant:6.93:DC;ADA2A::::6.9:C;5HT6R::::6.9:C;DRD1::BOVIN::6.89:C;DRD2:::ant:6.77:DC;5HT2B::::6.66:C;ACM2:::ant:6.41:DC;DRD5::RAT::5.98:C;ACM1::RAT::5.95:C;DRD1:::ant:5.91:DC;HRH1::RAT::5.9:C;HRH2::::5.55:C;5HT1A::RAT::5.53:C;HIF1A::::5.3:C;PRIO::::5.3:C;SCN1A::::5.27:C;P53::::5.:C;LEF::BACAN::5.:C;ADA1A:::ant::D;ADA1B:::ant::D;DRD4:::ant::D|CP2D6:::sub:7.3:DC;CP1A2:::inh:5.9:DC;CP2CJ:::sub:5.1:DC;CP2C9:::sub::D;CP3A4:::sub::D||
Spironolactone|ok|MCR:::ant:8.8:DC;GCR:::ant:7.49:DC;ANDR:::ant:7.4:DC;ANDR::RAT::7.04:C;PRGR:::ago:6.4:DC;CP2CJ::::5.52:C;ESR2::::5.48:C;ESR1::::5.24:C;NR1I2;CCG1,CCG2,CCG3,CCG4,CCG5,CCG6,CCG7,CCG8,CA2D1,CA2D2,CA2D3,CA2D4,CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1B,CAC1A,CAC1E,CAC1G,CAC1H,CAC1I:::inh::D;SHBG:::bin::D;S5A1,S5A2,PORED:::ant::D;CP17A:::ant::D;C11B2:::ant::D|C11B1:::ind::D;CP2C8:::inh::D|ABCBB:::sub::D;SO1A2:::inh::D;MDR1:::ind::D;MRP2:::ind::D|A1AG1,A1AG2;ALBU
Methylphenidate|ok_inv|SC6A3:::inh:7.77:DC;SC6A2:::inh:7.21:DC;SC6A3::RAT::7.08:C;SC6A4::::5.29:C;5HT1A|Q6LAP9:::sub::D||
Methocarbamol|ok_vet|CAH1:::inh::D|||
Hyoscyamine|ok|AMPC::ECOLI::5.05:C;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D|||
Zolpidem|ok|GBRA1:::ago:7.85:DC;GBRG2::RAT::7.72:C;GBRP::RAT::7.6:C;GBRG2:::ago:6.99:DC;GBRB2::::6.74:C;GBRA2:::ago:6.13:DC;GBRA2::RAT::6.12:C;TSPO::RAT::5.33:C;LMNA::::5.25:C;GBRA3:::ago::D|CP2D6:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP1A2:::sub::D;CP3A4:::sub::D||
Famciclovir|ok_inv|DPOL::VZVD:inh::D;DPOL::HHV11:inh::D|AOXA:::sub::D||
Triprolidine|ok|HRH1::CAVPO::9.9:C;HRH1:::ant:8.8:DC|||
Streptozocin|ok_inv|OGA;OGA::BACTN:ant::D;GTR2:::lig::D;DNA:::cov::D|CP2E1:::ind::D;CP1A2:::ind::D;CP1A1:::ind::D|MDR1:::ind::D|
Carboprost_tromethamine|ok|PE2R1:::ago::D|||
Cefpiramide|ok|PBP2A::STAAU:inh::D;PBPA::ECOLI:inh::D;DACC::ECOLI:inh::D;Penicillin_binding_protein_1B::PSEAI:inh::D;PBPA::PSEAE:inh::D;PBPB::ECOLI:inh::D;FTSI::ECOLI:inh::D|||ALBU
Lindane|ok_out|GBRB3::::9.05:DC;GBRG2::::8.31:C;GBRB::MUSDO::7.96:C;GBRA1::::7.68:C;GBRR1::::7.04:DC;NR1I2;ESR1;PRGR;GLRB:::ant::D;GLRA3:::ant::D;GLRA2:::ant::D;GLRA1:::ant::D;GBRB1:::ant::D|||
Trifluridine|ok_inv|LMP1::EBVB9::5.95:C;LMNA::::5.7:C;AMPC::ECOLI::5.25:C;DNA;TYSY:::inh::D|TYPH:::sub::D;KITH:::sub::D|S29A2:::sub::D;S29A1:::sub::D;S28A1:::sub::D;S22A6:::inh::D|ALBU:::bin::D
Prochlorperazine|ok_vet|5HT2A::::8.7:C;HRH1:::ant:8.55:DC;DRD2:::ant:8.44:DC;DRD3::::8.35:C;ADA2B::::8.32:C;ADA2C::::7.92:C;ADA1A::RAT::7.89:C;ADA1D::::7.8:C;SGMR1::::7.64:C;5HT2C::::7.39:C;ADA1B::RAT::7.31:C;ADA2A,ADA2B,ADA2C:::ant:7.2,8.32,7.92:DC;ADA2A::::7.2:C;5HT2B::::7.19:C;DRD1::::7.11:C;LMNA::::7.05:C;5HT6R::::6.91:C;ACM5::::6.8:C;ACM4::::6.72:C;5HT4R::CAVPO::6.71:C;ACM1::::6.61:C;ACM3::::6.49:C;SC6A2::::6.4:C;5HT1A::RAT::6.27:C;SC6A4::::6.21:C;DRD4::::6.09:C;CP1A2::::6.:C;ACM2::::5.96:C;5HT1B::RAT::5.92:C;SC6A3::::5.86:C;KCNH2::::5.82:C;PDR5::YEAST::5.77:C;CP2CJ::::5.7:C;TSHR::::5.5:C;MCL1::::5.42:C;CP3A4::::5.3:C;ACM1::RAT::5.25:C;FYN::::5.25:C;MK01::::5.:C;ADA1A,ADA1B,ADA1D:::ant:,,7.8:DC|CP2D6:::sub:6.52:DC||
Cyproheptadine|ok|5HT2A:::ant:9.56:DC;HRH1:::ant:9.37:DC;HRH1::CAVPO::9.27:C;5HT2C:::ant:8.89:DC;5HT2A::RAT::8.8:C;ACM4::::8.66:C;ACM5::::8.56:C;5HT2B::RAT::8.51:C;ACM1:::ant:8.4:DC;ACM1::RAT::8.4:C;5HT2B::::8.22:C;5HT3A::RAT::8.1:C;ACM3:::ant:8.02:DC;5HT2C::MOUSE::7.96:C;ACM2:::ant:7.92:DC;DRD3::::7.8:C;ADA2B::::7.77:C;ADA1B::RAT::7.36:C;5HT7R::::7.3:DC;5HT7R::RAT::7.3:C;ADA1D::::7.28:C;DRD2::::7.26:C;DRD5::RAT::7.2:C;5HT1A::RAT::7.15:C;DRD1::::7.1:C;ADA1A::RAT::7.01:C;ADA2A::::6.97:C;DRD2::MOUSE::6.95:C;5HT6R::::6.89:C;DRD2::RAT::6.85:C;ADA2C::::6.73:C;HRH2::::6.71:C;SC6A2::MOUSE::6.54:C;SC6A2::::6.54:C;TSHR::::6.:C;SETD7::::6.:C;SCN1A::::6.:C;5HT1B::RAT::5.9:C;CP2D6::::5.6:C;LEF::BACAN::5.4:C;SC6A4::MOUSE::5.39:C;SC6A4::::5.39:C;CAC1C::CAVPO::5.11:C|UD13:::sub::D||
Nitric_Oxide|ok|GCYA2:::ind::D;MT1A;I23O1|ALDH2:::inh::D;CP1A2:::inh::D;CP2B6:::inh::D;CP3A4:::inh::D||
Bendroflumethiazide|ok|LMNA::::6.3:C;CAH4:::inh::D;CAH2:::inh::D;CAH1:::inh::D;KCMA1:::ind::D;S12A3:::inh::D|TPMT:::inh::D||
Allopurinol|ok|XDH::BOVIN::6.59:C;BLM::::6.4:C;XDH::RAT::6.12:C;RAB9A::::6.:C;TSHR::::5.3:C;LMNA::::5.2:C|XDH:::inh:8.44:DC;AOXA:::sub::D|S22A2;ABCG2:::sub::D;S22A7:::sub::D;S22A8:::sub::D|
Ceftazidime|ok|PBP5::PSEAE:inh::D;MRDA::ECOLI:inh::D;Penicillin_binding_protein_2::PSEAI:inh::D;Penicillin_binding_protein_1B::PSEAI:inh::D;PBPB::ECOLI:inh::D;PBPA::STRR6:inh::D;PBPA::ECOLI:inh::D;PBP3::STREE:inh::D;FTSI::ECOLI:inh::D||S22A6:::inh::D;S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|
Cerivastatin|ok_out|HMDH:::inh:10.07:DC;HMDH::RAT::8.55:C|UD11:::sub::D;CP2B6:::ind::D;CP2C9:::inh::D;CP2D6:::inh::D;CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::duo::D|ABCBB:::sub::D;SO1B1:::inh::D;ABCG2:::sub::D;MRP2:::sub::D;MDR1:::sub::D|
Trimethoprim|ok_vet|DYR::STAAU::8.92:C;DYR::CANAX::8.66:C;BLM::::8.49:C;HCD2::::8.2:C;DRTS::TOXGO::8.14:C;DRTS::PLAFK::8.:C;DYR:::inh:8.:DC;DYR::PNECA::7.34:C;DYR::LACCA::7.27:C;DRTS::PLABA::6.92:C;DRTS:S108N:PLAFK::6.88:C;NFKB1::::6.6:C;DYR::LACLA::6.35:C;DYR::NEIGO::6.35:C;DYR1::ECOLX::6.3:C;DYR::MOUSE::6.3:C;DYR::ECOLI::5.57:C;TSHR::::5.3:C;TYSY:::inh::D|CP2C9:::sub::D;CP2C8:::inh::D;CP3A4:::sub::D|S22A2:::inh::D;MDR1:::duo::D|
Gemcitabine|ok|KCY:::inh::D;TYSY:::inh::D;RIR1:::inh::D;DNA:::cov::D|DCK:::sub::D;CDD:::sub::D|S28A3:::sub::D;S29A2;S28A1;S29A1:::sub::D;MRP7:::sub::D;MDR1:::sub::D|
Entecavir|ok_inv|DNA|||
Betamethasone|ok_vet|GCR:::ago:8.45:DC|CP3A5:::ind::D;CP19A:::sub_ind::D;CP3A4:::sub_ind::D|MDR1:::sub::D|
Teniposide|ok|TOP2A:::inh::D|CP3A5:::sub::D;CP2CJ:::sub::D;CP2C9:::inh::D;CP3A4:::inh::D|ABCG2:::sub::D;MRP6:::sub::D|
Epirubicin|ok|5HT4R::CAVPO::5.88:C;FYN::::5.29:C;DNA:::itc::D;TOP2A:::inh::D;CHD1:::ant::D|PA24A:::inh::D;UD2B7:::sub::D|MRP1:::sub::D|
Chloramphenicol|ok_vet|STRP::STRP1::6.01:C;DAF;DRAA::ECOLX:ant::D;RL16::ECOLI:inh::D|CPT::STRVP:sub::D;CAT4::PSEAE:sub::D;CAT3::ECOLX:sub::D;CP2CJ:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D|S22A6:::inh::D|
Loracarbef|ok_out|PBPA::CLOPE:inh::D;PBP3::STREE:inh::D||S15A2:::inh::D;S15A1:::inh::D|
Lansoprazole|ok_inv|TAU::::8.6:DC;ACM1::RAT::7.25:C;TSHR::::6.9:C;LMNA::::6.9:C;ATP4A:::inh:6.4:DC;PHOP1::::6.36:C;HCD2::::6.3:C;NPC1::::5.64:C;RAB9A::::5.64:C;AGAL::::5.3:C;FAS::::5.28:C;CP1A2::::5.19:C;HIF1A::::5.1:C;I23O2::MOUSE::5.09:C|CP2CJ:::inh:7.:DC;CP2D6:::inh:5.54:DC;CP2C8:::sub:5.24:DC;CP3A4:::duo::D;CP2CI:::sub::D;CP2C9:::duo::D;CP1B1:::ind::D;CP1A1:::ind::D|S22A3;S22A2;S22A1;S22A8:::inh::D;MDR1:::inh::D;ABCG2:::inh::D|
Dipivefrin|ok|ADA1A:::ago::D;ADA2A:::ago::D;ADRB2:::ago::D;CHLE:::sub::D;ACES:::inh::D|||
Droperidol|ok_vet|ADA1A::RAT::9.17:C;5HT2A::::9.13:C;DRD2:::ant:9.1:DC;DRD3::::9.03:C;ADA1B::RAT::8.01:C;KCNH2::::7.49:C;ADA1D::::7.39:C;ADA2B::::7.:C;5HT1A::RAT::6.86:C;5HT2C::::6.62:C;ADA2C::::6.59:C;HRH1::::6.28:C;ACM4::::6.27:C;DRD1::::6.26:C;5HT4R::CAVPO::6.2:C;SCN1A::::6.13:C;5HT2B::::6.07:C;ADA2A::::5.95:C;ACM5::::5.78:C;LEF::BACAN::5.6:C;CP2D6::::5.5:C;HIF1A::::5.4:C;MK01::::5.35:C;CP3A4::::5.2:C;CAC1C::::5.12:C;RORG::MOUSE::5.1:C;ADA1A:::ant::D|||
Levothyroxine|ok|LMNA::::6.15:C;NR1H4::::5.1:C;ITB3;ITAV;THB:::ago::D;THA:::ago::D|UD11:::sub:5.31:DC;CP2C8:::inh::D|SO4C1::::5.1:DC;SO2B1:::inh::D;LAT1;SO4A1;SO1B3:::inh::D;SO1B1:::inh::D;SO1A2:::inh::D;MOT8:::inh::D;SO1C1:::inh::D;MDR1:::ind::DC|TTHY::::5.66:DC;ALBU;THBG:::sub::D
Framycetin|ok|TRPV1::::6.4:C;LEF::BACAN::6.3:C;CXCR4:::ant::D;RS12::ECOLI:inh::D;16S_ribosomal_RNA::Gut_flora:inh::D|||
Clomocycline|exp|RS4::ECOLI:inh::D;RS9::ECOLI:inh::D;16S_ribosomal_RNA::Gut_flora:inh::D|||
Meperidine|ok|OPRM:::ago:6.5:DC;KCNH2::::6.49:C;SC6A4::RAT::6.39:C;OPRM::CAVPO::6.35:C;OPRK::::6.3:DC;OPRM::MOUSE::6.3:C;SGMR1::RAT::6.15:C;EST1;SC6A4:::bin::D;SC6A2:::inh::D;SC6A3:::inh::D;ACM1,ACM2,ACM3,ACM4,ACM5:::bin::D;NMDE4:::ant::D;NMDE3:::ant::D;NMDE1:::ant::D;NMDE2:::ant::D;NMDZ1:::ant::D|CP1A2:::ind::D;CP2D6:::sub::D;CP2B6:::sub::D;CP2CJ:::sub::D;CP3A4:::sub_ind::D||A1AG1;ALBU
Loratadine|ok_inv|HRH1:::ant:7.7:DC;HRH1::CAVPO::7.14:C;5HT2B::::6.81:C;KCNH2:::ant:6.77:DC;HRH1::RAT::6.46:C;ACM1::RAT::5.9:C;NR1I2::::5.52:C;NR1H4::::5.51:C;MEN1::::5.45:C;S6A15::::5.4:C;NPSR1::::5.4:C;TAU::::5.:C|CP2CJ:::inh:7.8:DC;CP2C9:::sub:7.4:DC;CP2C8:::inh:5.53:DC;CP3A4:::inh:5.2:DC;UDB15;UD13;UD11;UDB10;CP3A5:::sub::D;CP2B6:::sub::D;CP1A2:::sub::D;CP1A1:::sub::D;CP2D6:::inh::D|ABCBB:::sub::D;MDR1:::inh::D|
Cefalotin|ok_inv_vet|CTDS1::::5.56:C;DNMT1::::5.14:C;AMPC::ECOLI:pot::D;PBPA::CLOPE:inh::D;PBP2::STRR6:inh::D;PBP2A::STRR6:inh::D;PBP3::STREE:inh::D;PBP1B::STRR6:inh::D;PBPA::STRR6:inh::D;DAC::STRSR:inh::D||S22A8:::inh:7.4:DC;S22AB:::inh:6.7:DC;S22A6:::inh:6.66:DC;S22A7:::inh::D;S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|ALBU:::bin::D
Prazosin|ok|ADA1B::RAT::10.99:C;ADA1A,ADA1B,ADA1D::::10.4,9.68,9.7:DC;ADA1A:::ant:10.4:DC;ADA1A::RAT::10.15:C;ADA1A::BOVIN::9.9:C;ADA1D::RAT::9.77:C;ADA1D:::ant:9.7:DC;OPRM::RAT::9.7:C;ADA1B:::ant:9.68:DC;5HT1D::::9.48:C;CASB::RAT::9.44:C;ADA2C::RAT::9.4:C;ADA1B::MESAU::9.16:C;AA3R::::9.07:C;ADA1A::RABIT::8.3:C;ADA2B::RAT::8.11:C;NQO2::::8.11:C;ADA2B:::bin:7.89:DC;ADA2B::MOUSE::7.89:C;ADA2C::::7.62:C;ADA2A:::bin:7.47:DC;ADA2A::BOVIN::6.97:C;LMNA::::6.95:C;KDM4E::::6.2:C;5HT2A::RAT::5.82:C;KCNH2:::inh:5.8:DC;S47A1::::5.8:C;ADA2A::RAT::5.78:C;5HT1A::RAT::5.63:C;5HT2B::::5.58:C;SMN::::5.4:C;MMP1::::5.39:C;ADA2A::PIG::5.39:C;HD::::5.35:C;CP3A4::::5.2:C;MMP9::::5.16:C;LEF::BACAN::5.1:C;DRD4::::5.08:C;SCN1A::::5.:C||S22A1:::inh:5.74:DC;ABCG2:::sub::D;MDR1:::inh::D;S22A3:::inh::D|A1AG1:::sub::D
Imipramine|ok|HRH1::RAT::10.22:C;SC6A4:::inh:9.28:DC;ADA1A::RAT::8.77:C;SC6A4:W103A::inh:8.59:DC;AA3R::::8.36:C;SC6A4::MOUSE::8.3:C;SC6A4:I179C::inh:8.24:DC;SC6A2::MOUSE::7.92:C;SC6A2:::inh:7.8:DC;5HT2B::RAT::7.64:C;HRH1:::ant:7.57:DC;SC6A3::MOUSE::7.38:C;SC6A4::RAT::7.38:C;5HT3A::RAT::7.36:C;ADA1B::RAT::7.34:C;ACM1::RAT::7.19:C;5HT2A:::ant:7.03:DC;5HT2C::MOUSE::6.8:C;5HT2C:::ant:6.8:DC;ADA2C::RAT::6.59:C;ACM5::RAT::6.52:C;DRD2:::bin:6.39:DC;TAU::::6.25:C;DRD5::RAT::6.19:C;DRD2::MOUSE::6.14:C;LMNA::::6.1:C;SC6A4:I172M::inh:5.89:DC;HRH2::CAVPO::5.72:C;KCNH2:::inh:5.47:DC;SCN1A::::5.44:C;CAC1C::RAT::5.39:C;MTOR::::5.28:C;AL1A1::::5.25:C;CAC1C::::5.08:C;S22A2::RAT::5.:C;PRIO::::5.:C;S47A1::::5.:C;A1AG2;KCNH1;5HT6R:::bin::D;5HT1A:::act::D;SC6A3:::inh::D;DRD1,DRD5:::bin::D;5HT7R:::ant::D;ADA1B:::ant::D;KCND3:::inh::D;KCND2:::inh::D;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;ADA1D:::ant::D;ADA1A:::ant::D|CP2D6:::inh:5.2:DC;CP2E1:::inh::D;CP2CI:::sub::D;CP2B6:::sub::D;CP3A7:::sub::D;CP3A4:::sub::D;CP1A2:::inh::D;CP2CJ:::inh::D|S22A2:::inh:6.22:DC;S22A4:::inh::D;S22A3:::inh::D;MDR1:::sub::D|ALBU;A1AG1
Acitretin|ok|SMN::::5.5:C;RET1:::ago::D;RXRG:::ago::D;RXRB:::ago::D;RARG:::ago::D;RARB:::ago::D;RARA:::ago::D;RXRA:::ago::D|||ALBU
Verteporfin|ok_inv||||
Nabumetone|ok|LMNA::::6.25:C;AOFA::::6.:C;SC6A2::::5.73:C;NPC1::::5.55:C;RAB9A::::5.55:C;KDM4E::::5.15:C;PGH1:::inh::D;PGH2:::inh::D|CP1A2:::sub:6.4:DC;AK1C4:::sub::D;AK1C2:::sub::D;AK1C1:::sub::D;DHI1:::sub::D;CP2C9:::sub::D;PERM:::inh::D||ALBU
Methscopolamine_bromide|ok|ACM1:::ant::D;ACM2:::ant::D;ACM3:::ant::D|||
Metharbital|out|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA4:::pot::D;GBRA5:::pot::D;GBRA6:::pot::D;ACHA4:::ant::D;ACHA7:::ant::D;GRIA2:::ant::D;GRIK2:::ant::D;GABAR:::aga::D|||
Sodium_tetradecyl_sulfate|ok_inv|PROS:::inh::D;PROC:::inh::D|||
Ketorolac|ok|PGH1:::inh:7.89:DC;PTGDS::MOUSE::6.64:C;PGH2:::inh:6.37:DC;RAB9A::::5.44:C;ALDR::RAT::5.21:C|CP2C9:::sub::D;CP2C8:::sub::D;UD2B7:::sub::D||
Enoxacin|ok_inv|LMNA::::5.9:C;VATB2::::5.:C;TOP2A:::inh::D;PARC::HAEIN:inh::D;GYRA::HAEIN:inh::D|CP1A2:::inh::D||
Quinine|ok|S22A1::MOUSE::6.55:C;S22A1::RAT::6.05:C;S22A2::MOUSE::5.55:C;SO1A4::RAT::5.42:C;SCN1A::::5.36:C;KCNN4:::inh::D;GPIX;Fe_II_protoporphyrin_IX::PLAFA:ant::D|CP2D6:::inh:5.74:DC;CP3A4:::duo::D;CP1A1:::duo::D;CP3A7:::sub::D;CP2E1:::sub::D;CP2CJ:::inh::D;CP2C9:::sub::D;CP2C8:::inh::D;CP1A2:::sub::D;CP3A5:::sub::D|S22A2:::inh:5.47:DC;SO1B1:::inh::D;S22A4:::inh::D;SO1A2:::inh::D;MDR1:::inh::D;S22A5:::inh::D;S22A1:::inh::D|
Tenoxicam|ok|LYAG::::6.:C;PGH1:::inh:5.94:DC;KDM4E::::5.05:C;PGH2:::inh::D|CP2C9:::sub:5.6:DC|S22A8:::inh::D|
Dronabinol|ok_ill|CNR2:::ago:8.82:DC;CNR1:::ago:8.55:DC;CNR2::RAT::8.24:C;CNR1::RAT::8.24:C;CNR2::MOUSE::8.04:C;CNR1::MOUSE::7.82:C;TRPA1::RAT::6.64:C;GPR18::::6.02:C;GLRA1::::5.89:C|PGH1:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D|ABCG2:::inh::D;MDR1:::inh::D|
Montelukast|ok|CLTR1:::ant:9.37:DC;CLTR1::CAVPO::9.3:C;AA3R::::6.61:C;ADA2C::::6.12:C;MK14::::6.07:C;NK2R::::5.89:C;ACM3::::5.85:C;ADA2A::::5.83:C;THAS::::5.82:C;OPRD::::5.77:C;ACM1::::5.71:C;SC6A3::::5.68:C;ADRB2::::5.62:C;DRD3::::5.58:C;SC6A2::::5.57:C;EGFR::::5.5:C;ADRB3::::5.49:C;5HT2B::::5.4:C;FYN::::5.33:C;GPR17::::5.18:C;LOX5|CP2A6:::sub::D;PGH1:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D;CP2C8:::inh::D|SO2B1:::sub::D|
Fluoxetine|ok_vet|SC6A4:::inh:9.57:DC;SC6A4::RAT::8.57:C;ADA2A::::8.2:C;KCNH2:::inh:8.:DC;SC6A3::MOUSE::7.97:C;5HT1B::RAT::7.82:C;5HT2A::::7.26:C;5HT2C:::ant:7.21:DC;SC6A2::MOUSE::7.07:C;5HT2C::RAT::6.96:C;ACES::::6.89:C;SGMR1::::6.68:C;SC6A2::::6.62:C;ADA1B::RAT::6.22:C;ADA2B::::6.16:C;ACM3::::6.12:C;ACM1::::6.11:C;5HT6R::::6.11:C;ACM5::::6.01:C;SC6A3::RAT::5.96:C;LMNA::::5.85:C;ADA2C::RAT::5.72:C;SC6A3::::5.72:C;CAC1C::RAT::5.55:C;CAC1C::::5.27:C;HRH3::::5.14:C;CKS1;ACHB4:::ant::D;ACHA3:::ant::D;ACHA2:::ant::D|CP2CJ:::inh:7.4:DC;CP2D6:::inh:6.15:DC;CP3A5:::sub::D;CP2B6:::sub::D;CP3A4:::inh::D;CP1A2:::inh::D;Q14097:::ind::D;CP2C9:::inh::D|MDR1:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Hexylcaine|ok_out|SCN1A::::5.15:C;SCNAA:::inh::D;SCN5A:::inh::D|||
Methohexital|ok|GBRA1:::ant::D|CP2CJ:::sub::D||
Chlordiazepoxide|ok_ill_inv|GBRP::RAT::6.7:C;HRH1::::6.68:C;GBRG2::::6.56:C;TSPO::RAT::6.36:C;GBRA1::::6.25:C;GBRA2::BOVIN::6.1:C;GABAR:::aga::D|||
Duloxetine|ok|SC6A4::RAT::10.09:C;SC6A4:::inh:9.62:DC;SC6A2:::inh:8.8:DC;SC6A3:::inh:6.62:DC;SC6A3::RAT::6.43:C;CP3A4::::6.36:C;CAC1C::::5.55:C;CP2CJ::::5.39:C;KCNH2::::5.3:C;KMT2A::::5.15:C;SCN5A::::5.1:C;KCNQ1::::5.:C|CP2D6:::inh:6.:DC;CP1A2:::sub:5.28:DC;CP2C9:::sub::D|MDR1:::inh::D|A1AG1,A1AG2:::lig::D;ALBU:::lig::D
Chlorpromazine|ok_inv_vet|5HT2B::RAT::9.15:C;DRD2:::ant:9.:DC;5HT2A,5HT2B,5HT2C:::bin:8.96,7.4,8.56:DC;5HT2A:::ant:8.96:DC;DRD2::RAT::8.92:C;DRD3:::inh:8.8:DC;ADA1B::RAT::8.8:C;HRH1:::ant:8.71:DC;ADA1D::::8.71:C;DRD1::RAT::8.67:C;5HT2C:::bin:8.56:DC;ADA1A::RAT::8.46:C;5HT6R:::bin:8.4:DC;DRD5::RAT::8.01:C;5HT7R:::bin:7.97:DC;ADA2B::::7.92:C;ACM5::::7.74:C;SC6A2::::7.72:C;ACM1:::ant:7.7:DC;ACM4::::7.68:C;SC6A4::::7.68:C;5HT7R::RAT::7.68:C;DRD4:::bin:7.6:DC;DRD1::BOVIN::7.6:C;5HT2B::::7.4:C;ACM3:::ant:7.36:DC;HRH1::CAVPO::7.3:C;ADA2C::::7.27:C;ACM1::RAT::7.22:C;DRD2::BOVIN::7.1:C;DRD1,DRD5:::inh:7.02,6.76:DC;DRD1:::ant:7.02:DC;ADA2A,ADA2B,ADA2C:::inh:6.88,7.92,7.27:DC;ADA2A::::6.88:C;DRD5:::inh:6.76:DC;5HT1A::RAT::6.75:C;SGMR1::::6.72:C;LMNA::::6.65:C;ACM2::::6.63:C;ADA2C::RAT::6.3:C;TRPV1::RAT::6.28:C;AOXA::::6.24:C;NMDZ1::::6.22:C;5HT1A:::ant:6.17:DC;CALM1:::inh:5.91:DC;ACHA::TETCF::5.89:C;NMDZ1::RAT::5.89:C;KCNH2:::inh:5.83:DC;5HT1B::RAT::5.74:C;PRIO::::5.7:C;SC6A3::::5.68:C;CALM::BOVIN::5.6:C;HRH2::::5.59:C;KCNK2::::5.57:C;TYTR::TRYCR::5.49:C;CAC1C::::5.47:C;SCN1A::::5.37:C;S22A1::::5.37:C;PDR5::YEAST::5.35:C;OPRK::::5.35:C;OPRM::::5.23:C;MC5R::::5.15:C;OPRD::::5.13:C;FYN::::5.06:C;NK2R::::5.04:C;P53::::5.:C;LEF::BACAN::5.:C;HRH4:::bin::D;A1AG1,A1AG2:::bin::D;ASM:::inh::D;ADA1A,ADA1B,ADA1D:::inh:,,8.71:DC;ADA1B:::ant::D;ADA1A:::ant::D|CP2D6:::inh:6.8:DC;CP3A4:::ind:6.:DC;CP1A2:::sub:6.:DC;CHLE:::inh::D;CP2E1:::inh::D|MDR1:::inh:6.22:DC;ABCBB:::inh::D|ALBU
Rimantadine|ok_inv|M2::I000F::7.8:C;S22A2::::5.36:C;S47A1::::5.14:C;M2::I60A0:::D|||
Amikacin|ok_inv_vet|LMNA::::6.8:C;RS12::ECOLI:inh::D|||
Lenalidomide|ok|PGH2:::neg::D;CADH5:::ant::D;TNF11:::inh::D;CRBN:::inh::D||MDR1:::sub::D|
Raloxifene|ok_inv|ESR1:::ago:10.52:DC;ESR2:::ago:9.7:DC;ESR1::RAT::9.15:C;EBP::::9.:C;ESR2::RAT::8.47:C;SGMR1::::7.42:C;ERG2::YEAST::7.18:C;5HT2B::::7.16:C;ADA2C::::6.97:C;SC6A2::::6.55:C;LMNA::::6.45:C;DRD2::::6.41:C;ACES::::6.4:C;5HT2A::::6.38:C;OPRM::::6.32:C;ADA1D::::6.32:C;AOXA::MOUSE::6.3:C;AOXA::MACFA::6.3:C;AL1A1::::6.3:C;DRD3::::6.27:C;5HT2C::::6.21:C;ADA2A::::6.2:C;OPRK::::6.19:C;5HT6R::::6.12:C;5HT1B::RAT::6.07:C;ADA1A::RAT::6.05:C;AOXA::RAT::5.96:C;AA2AR::::5.93:C;NK2R::::5.88:C;ADA1B::RAT::5.83:C;SC6A3::::5.83:C;ADA2B::::5.77:C;SC6A4::::5.72:C;DRD1::::5.71:C;CP2C9::::5.7:C;OPRD::::5.63:C;HCD2::::5.6:C;PLD2::::5.47:C;FYN::::5.44:C;PLD1::::5.4:C;LEF::BACAN::5.3:C;CP2CJ::::5.2:C;CP2D6::::5.1:C;TFF1;SPB9|AOXA:::inh:9.06:DC;CP3A4:::inh:5.9:DC;UD18:::sub::D;UD110:::sub::D;UD11:::sub::D;CP19A:::inh::D;CP2C8:::inh::D;CP2B6:::inh::D|MRP4:::sub::D;MRP3:::sub::D;MRP2:::sub::D;ABCG2:::sub::D;MDR1:::sub::D;SO1B3:::sub::D;SO1B1:::sub::D|A1AG1:::bin::D;ALBU:::bin::D
Celecoxib|ok_inv|PGH2::MOUSE::9.29:C;PGH2:::inh:9.28:DC;PGH1::MOUSE::9.15:C;PGH1::SHEEP::8.43:C;CAH9::::7.8:C;CAH12::::7.74:C;CAH2:::inh:7.68:DC;CAN::CANAL::7.68:C;PGH2::SHEEP::7.4:C;CAH15::MOUSE::7.35:C;PGH1::::7.3:C;PGH2::BOVIN::7.24:C;COX2::SHEEP::7.22:C;CAH6::::7.03:C;CAH5B::::7.03:C;CAH13::::7.01:C;CAN::YEAST::6.97:C;CAH::METTE::6.85:C;PGH2::RAT::6.85:C;CAH4::BOVIN::6.54:C;PTGES::::6.37:C;ADA2B::::6.16:C;CAH14::::6.16:C;MTCA2::MYCTU::6.15:C;CAH5A::::6.1:C;TSHR::::6.1:C;MK14::::6.09:C;CAH4::::6.06:C;SC6A3::::5.71:C;CAH7::::5.66:C;SC6A4::::5.48:C;PGH1::CANLF::5.25:C;SC6A2::::5.14:C;CAH3:::inh:5.13:DC;PGH1::BOVIN::5.11:C;Cadherin_11:::inh::D;PDPK1:::inh::D|CP2D6:::inh:6.:DC;CP2C9:::sub:5.:DC;CP2C8:::sub::D;CP3A4:::sub::D|ABCG2:::sub::D;MDR1:::sub::D;ABCBB:::inh::D;MRP4:::inh::D|
Gallamine_triethiodide|ok|ACM2:::ant:6.15:DC;ACM5;ACM1;ACHA2:::ant::D;ACES:::inh::D|||
Brimonidine|ok|ADA2A:::ago:9.21:DC;ADA2C:::ago:8.47:DC;ADA2C::RAT::8.44:C;BLM::::8.25:C;ADA2B:::ago:7.46:DC;ADA2B::RAT::7.28:C;CP3A4::::6.4:C;ADA1B::RAT::6.13:C;ADA1D::::6.07:C;ADA1A::::5.96:C;ADA1A::BOVIN::5.95:C;5HT1A::RAT::5.84:C;LMNA::::5.6:C;ADA1A::RAT::5.59:C;KDM4E::::5.45:C;ADA1B::::5.36:C;END4::ECOLI::5.1:C|AOXA:::sub::D||
Dicloxacillin|ok_inv_vet|PBP2::STRR6:inh::D;PBPA::STRR6:inh::D;PBP2A::STRR6:inh::D;PBP1B::STRR6:inh::D;PBP3::LISMN:inh::DC|CP3A4:::ind::D|S15A2:::inh::D;S15A1:::inh::D|
Nabilone|ok_inv|CNR2:::pag:8.74:DC;CNR2::MOUSE::8.74:C;CNR1:::pag:8.66:DC;CNR1::RAT::8.66:C|CP2C9:::inh::D;CP2C8:::inh::D;CP2E1:::inh::D||
Pefloxacin|ok|TOP1::STAAU:inh::D;TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A2:::inh::D||
Altretamine|ok|THB::::8.8:C;HCD2::::6.5:C;LMNA::::6.1:C;CP1A2::::5.7:C;ACM1::RAT::5.55:C;DNA|||
Sotalol|ok|LMNA::::8.46:C;ADRB2:::ant:6.53:DC;ADRB2::BOVIN::6.24:C;ADRB1:::ant:6.08:DC;ADRB2::CANLF::5.3:C;KCNH2:::inh::D|CP2D6:::sub::D||
Buspirone|ok_inv|5HT1A:::pag:8.51:DC;5HT1A::RAT::8.42:C;DRD2:::ant:7.89:DC;DRD3:::ant:7.82:DC;5HT1B::RAT::7.77:C;SGMR1::::7.44:C;DRD2::RAT::7.38:C;DRD2::BOVIN::7.36:C;SGMR1::RAT::7.32:C;DRD5::RAT::6.92:C;ADA1B::RAT::6.86:C;5HT2B::RAT::6.76:C;5HT2A::BOVIN::6.75:C;5HT2A::RAT::6.32:C;5HT2B::::6.32:C;ADA1D::::6.28:C;ADA1A,ADA1B,ADA1D:::pag:6.24,,6.28:DC;ADA1A::::6.24:C;5HT2A::::6.19:C;5HT2C::RAT::6.:C;ADA1A::RAT::5.85:C;S47A1::::5.77:C;5HT2C::::5.64:C;KCNH2::::5.4:C;AL1A1::::5.35:C;DRD1::BOVIN::5.21:C;CP2C9::::5.1:C;ADA2A::BOVIN::5.:C;ADA2C::RAT::5.:C;DRD4:::ant::D|CP2D6:::sub:5.:DC;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|A1AG1:::bin::D;ALBU:::bin::D
Miglitol|ok|SUIS::RAT::6.96:C;LYAG:::ant:6.46:DC;GDE::RABIT::6.41:C;LYAG::RAT::6.34:C;SUIS::::6.3:C;MGA:::ant:6.:DC;GANC:::ant::D;GANAB:::ant::D|AMYP:::inh::D||
Fosinopril|ok|ACE:::inh:9.:DC||S15A2:::sub::D;S15A1:::sub::D|
Cefotaxime|ok|Beta_lactamase::ACIBA:::D;ALBU;PBP2::STRR6:inh::D;PBPA::STRR6:inh::D;PBPC::BACSU:inh::D;PBP2A::STRR6:inh::D;PBP1B::STRR6:inh::D||S22A8:::inh:6.54:DC;S22A6:::inh:5.5:DC;S22AB:::inh:5.21:DC;S15A2:::inh::DC;S15A1:::inh::DC;S22A7:::inh::DC|
Entacapone|ok_inv|COMT::RAT::7.89:C;LMNA::::7.35:C;GPR35::::5.25:C|COMT:::inh:6.41:DC;CP2D6:::inh::D;UD19:::sub::D||
Zidovudine|ok|CXCR4::::8.1:C;TERT:::inh::D;Reverse_transcriptase_RNaseH::9HIV1:inh::D|KITH:::sub:5.54:DC;UD11:::sub_ind::D;UD2B7:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D;CP2A6:::sub::D|ABCG2:::sub::D;MRP5:::sub::D;MRP4:::sub::D;MDR1:::sub::D;S29A2;S28A1;S22AB;S22A8:::inh::D;S22A7;S22A6:::sub::D;S22A2|ALBU
Darifenacin|ok_inv|ADRB2::::9.1:C;ACM3:::ant:9.08:DC;ADRB2::CAVPO::9.:C;ACM5:::ant:8.64:DC;ACM3::RAT::8.6:C;ACM1:::ant:8.26:DC;ACM4:::ant:8.07:DC;ACM2:::ant:7.8:DC;ADRB1::::7.4:C;ACM2::RAT::7.2:C;KCNH2::::7.1:C;SCN5A::::5.8:C;ADRB1::RAT::5.64:C|CP2D6:::inh::D;CP3A4:::sub::D||
Oxycodone|ok_ill_inv|OPRM::RAT::7.36:C;OPRM::MOUSE::6.8:C;OPRM:::ago:6.3:DC;OPRD::RAT::5.96:C;OPRK::RAT::5.58:C;OPRD:::ago:5.4:DC;OPRK:::ago::D|CP3A5:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D||A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Phenindione|ok_inv|LMNA::::5.45:C;MK01::::5.25:C;P53::::5.:C;VKOR1:::inh::D|||
Flutamide|ok_inv|LMNA::::7.1:C;ANDR:::ant:6.81:DC;AAAD::::6.22:C;AMPC::ECOLI::6.2:C;END4::ECOLI::6.05:C;5HT4R::CAVPO::5.65:C;EST2::::5.64:C;ACM1::RAT::5.2:C;5HT6R::::5.08:C;ANDR::RAT::5.05:C;NR1I2;AHR:::ago::D|CP1A2:::sub:6.5:DC;CP3A4:::sub:5.3:DC;CP2CJ:::sub:5.:DC;CP3A5:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D||
Tolmetin|ok|PGH1:::inh:7.39:DC;IL8::::7.05:C;ALDR::RAT::5.67:C;ALDR::::5.62:C;PGH2:::inh::D|PERM:::inh::D;T23O:::inh::D|S22A6:::inh::D|ALBU
Cimetidine|ok_inv|HRH2:::ant:7.15:DC;ACM1::RAT::7.05:C;HRH2::RAT::6.6:C;HRH2::CAVPO::6.58:C;S22A1::MOUSE::6.23:C;ATP4A::::6.09:C;TSHR::::5.8:C;LMNA::::5.3:C;S22A1::RAT::5.24:C;MEN1::::5.2:C;S22A2::MOUSE::5.1:C;S22A2::RAT::5.03:C|FMO1:::sub::D;FMO3:::sub::D;CP2E1:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;C11B1:::inh::D;CP2D6:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D;CP2CJ:::inh::D;CP1A2:::inh::D|S47A1:::inh:5.92:DC;S47A2:::inh::D;ABCBB:::inh::D;S22A7:::inh::D;S22AB:::inh::D;S22A4:::inh::D;S22A8:::inh::D;S22A6:::inh::D;S22A5:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D;MDR1:::sub_ind::D|
Haloperidol|ok|DRD3:::ANT:10.22:DC;DRD2::RAT::10.12:C;DRD2:::ant:9.92:DC;SGMR1::::9.7:DC;DRD5::RAT::9.55:C;DRD2::BOVIN::9.52:C;ERG2::YEAST::9.3:C;SGMR1::RAT::9.19:C;DRD4::::9.13:C;SGMR1::CAVPO::9.08:C;ADA1B::RAT::9.:C;DRD1::BOVIN::8.74:C;DRD3::RAT::8.62:C;DRD3::CHLAE::8.52:C;5HT2B::RAT::8.38:C;DRD2::CHLAE::8.32:C;ADA1A::::8.24:DC;DRD1:::ant:8.21:DC;DRD1::PIG::8.02:C;KCNH2::::8.:C;DRD4::RAT::8.:C;5HT2B::::7.8:C;ADA1A::RAT::7.76:C;5HT2A::RAT::7.7:C;ADA1A::BOVIN::7.7:C;DRD1::RAT::7.7:C;5HT2A::::7.68:DC;AP2S1::RAT::7.62:C;5HT2B::MOUSE::7.58:C;5HT2A::BOVIN::7.52:C;5HT2A::PIG::7.52:C;DRD5::::7.42:C;ADA1D::::7.39:C;ACM1::RAT::7.27:C;EBP::::6.72:C;ACM2::RAT::6.62:C;5HT7R::RAT::6.58:C;ADA2C::::6.57:DC;NFKB1::::6.55:C;5HT7R::::6.5:DC;HRH1::::6.49:DC;HRH1::RAT::6.42:C;HRH1::CAVPO::6.4:C;5HT1A::RAT::6.4:C;ADA2B::::6.21:DC;H10::::6.11:C;OPRM::::6.:C;HRH2::::5.94:C;SCN1A::::5.92:C;CAC1C::::5.89:C;5HT1A::::5.82:DC;ACM1::::5.8:C;5HT2C::::5.76:DC;SC6A4::::5.74:C;SC6A2::::5.74:C;ADA2A::::5.73:DC;ADA2C::RAT::5.57:C;ACM5::::5.55:C;CP2J2::::5.33:C;5HT2C::RAT::5.33:C;ACM3::::5.33:DC;KCNK2::::5.26:C;5HT6R::::5.22:DC;TPO::::5.2:C;LEF::BACAN::5.:C;VMAT2;MCHR1;NMDE2:::ant::D|CP2CJ:::sub:5.54:DC;CP3A4:::inh:5.5:DC;CP2D6:::inh:5.44:DC;CP1A1:::sub::D;CP2C9:::sub::D;UD19:::sub::D;CBR1:::sub::D;CP1A2:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|MDR1:::inh:6.7:DC|
Ritonavir|ok_inv|THAS::::7.12:C;S47A1::::7.1:C;NK2R::::6.06:C;NR1I2:::act:5.4:DC;MK01::::5.4:C;SO1B3::::5.4:C;S47A2::::5.36:C;V1AR::::5.3:C;OPRK::::5.26:C;Pol_polyprotein::9HIV1:inh::D|CP2C9:::ind:7.8:DC;CP3A4:::duo:7.8:DC;CP3A5:::duo:6.92:DC;UD11:::ind:5.77:DC;CP2B6:::duo:5.7:DC;CP2D6:::inh:5.64:DC;CP343:::duo::D;CP3A7:::duo::D;CP2E1:::inh::D;CP1A2:::duo::D;CP2C8:::duo::D;CP2CJ:::duo::D|SO1B1:::inh:6.15:DC;MDR1:::duo:5.82:DC;SO2B1:::inh:5.23:DC;ABCBB:::sub::D;ABCG2:::inh::D;MRP2:::sub_ind::D;SO1A2:::inh::D;MRP1:::duo::D|ALBU
Levallorphan|ok|OPRM:::pag:9.32:DC;SGMR1::RAT::9.27:C;OPRM::RAT::9.2:C;OPRK::::9.17:C|||
Tridihexethyl|out|ACM3:::ant::D;ACM1:::ant::D;ACM2:::ant::D|||
Nitazoxanide|ok_inv_vet|RAB9A::::6.3:C;NPC1::::6.3:C;LEF::BACAN::5.9:C;RORG::MOUSE::5.55:C;NPSR1::::5.5:C;TSHR::::5.3:C;CP3A4::::5.1:C;ALDR::::5.09:C;LMNA::::5.05:C;P53::::5.:C|PFOR::DESAF:inh::DC||S19A1
Triflupromazine|ok_vet|ACM1::RAT::6.8:C;CP2D6::::6.4:C;CP1A2::::6.1:C;PDR5::YEAST::5.31:C;CHLE::HORSE::5.13:C;LEF::BACAN::5.:C;ACM2:::ant::D;ACM1:::ant::D;5HT2B:::ant::D;DRD2:::ant::D;DRD1:::ant::D|CHLE:::inh::D|MDR1:::inh::D|
Dextrothyroxine|ok_inv|THB:::ago:8.25:DC;THB::RAT::7.46:C;LMNA::::7.05:C;SO1C1::MOUSE::6.57:C;NMDZ1::RAT::6.48:C;CP2C9::::5.2:C;TTHY::::5.14:C;PERT;THA:::ago::D||LAT1;SO4C1;SO4A1;SO1C1;SO1B1|
Acetyldigitoxin|ok|AT1A1:::inh::D|||
Vancomycin|ok|SC6A4::RAT::7.3:C;ADA2A::::7.3:C;ADA2C::RAT::6.9:C;ADA1B::RAT::6.:C;MRAY::ECOLI::5.05:C;MURG::ECOLI::5.:C;D::G+Bac:lig::D|||HRH1::MOUSE:sub::D;A1AG1,A1AG2:::sub::D;ALBU:::sub::D
Aminocaproic_acid|ok_inv|THB::::6.4:C;LMNA::::5.9:C;RECQ1::::5.2:C;APOA;TPA:::ant::D;PLMN:::inh::D|AOXA:::sub::D||
Dextromethorphan|ok|SC6A4:::inh:8.84:DC;TSHR::::8.2:C;SGMR1::CAVPO::7.82:C;SGMR1:::ago:6.46:DC;SCN2A::RAT::5.89:C;NMDZ1::RAT::5.88:C;NMDZ1::::5.77:C;ACM1::RAT::5.4:C;SGMR1::RAT::5.29:C;CP2DQ::RAT::5.25:C;SC6A2:::inh::D;CY24B,CY24A,NCF1,NCF2,NCF4,RAC1,RAC2:::inh::D;OPRK:::ago::D;OPRD:::ago::D;OPRM:::ago::D;ACHA7:::ant::D;ACHB2:::ant::D;ACHB4:::ant::D;ACHA4:::ant::D;ACHA3:::ant::D;PGRC1:::bin::D;NMD3A:::ant::D;ACHA2:::ant::D;HCG20471_isoform_CRA_c:::ago::D|CP2D6:::sub:5.74:DC;CP2C9:::sub::D;CP2CJ:::sub::D;CP2B6:::sub::D;CP3A7:::sub::D;CP3A4:::sub::D||
Cisplatin|ok|DNA:::cov::D;3MG;A2MG;TRFE;ATOX1|PERM:::ind::D;XDH:::ind::D;CP4AB:::ind::D;PGH2:::inh::D;NAT::MYCTU:inh::D;CP2C9:::inh::D;CP2B6:::inh::D;CHLE:::inh::D;GSTT1:::sub::D;MT1A:::sub::D;MT2:::sub::D;SODC:::sub::D;GSTP1:::sub::D;NQO1:::sub::D;GSTM1:::sub::D|MRP3:::ind::D;MRP5:::ind::D;MRP2:::ind::D;S22A2:::inh::D;COPT1:::sub::D;COPT2:::sub::D;MRP6:::sub::D;MDR1:::sub::D;ATP7B:::sub::D;ATP7A:::sub::D;ABCG2:::sub::D|ALBU
Bentoquatam|ok||||
Anisotropine_methylbromide|ok|ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D|||
Albendazole|ok_vet|LMNA::::6.4:C;SMN::::5.3:C;PGDH::::5.2:C;FRDA::SHEON:inh::D;TBB4B:::inh::D;Tubulin_beta_2_chain::ASCSU:inh::D;TBA1A:::inh::D|CP1A2:::ind:6.4:DC;CP2CJ:::sub::D;CP3A4:::sub::D;CP1A1:::ind::D||
Trandolapril|ok|ACE:::inh:9.03:DC|EST1:::sub::D|S15A2:::sub::D;S15A1:::sub::D|
Caspofungin|ok|FKS1::ASPNC:inh::D|CP3A4:::inh::D|SO1B3:::sub::D;SO1B1:::inh::D;S22A6:::inh::D;MDR1:::inh::D;S22A1|
Carteolol|ok|ADRB1:::pag:8.72:DC;ADRB2:::ant::D|CP2D6:::sub::D||
Bentiromide|inv_out|HEPS:::lig::D|||
Alitretinoin|ok_inv|RARB:::ago:9.3:DC;RARG:::ago:9.1:DC;RXRA:::ago:8.82:DC;RXRB:::ago:8.59:DC;RXRG:::ago:8.4:DC;RXRG::MOUSE::8.4:C;RARA::MOUSE::8.15:C;RARB::MOUSE::8.15:C;RARA:::ago:8.15:DC;RXRB::MOUSE::7.92:C;RARG::MOUSE::7.77:C;RXRA::MOUSE::7.49:C;RXRA::RAT::6.96:C;RORG::MOUSE::5.1:C;CP26C;PSG5;IBP3||MDR1:::sub::D|RABP1:::ago::D;RABP2:::ago::D
Metolazone|ok|CAH7::::8.68:C;PGDH::::5.05:C;S12A3:::inh::D|||
Tolnaftate|ok_inv_vet|CP2CJ::::7.:C;CP2C9::::5.9:C;5HT2B::::5.89:C;CP1A2::::5.6:C;CP3A4::::5.4:C;LEF::BACAN::5.3:C;ERG1::CANAL:inh::D|||
Oxaliplatin|ok_inv|DNA:::cov::D|GSTT1:::sub::D;MT1A:::sub::D;MT2:::sub::D;PERM:::sub::D;SODC:::sub::D;GSTP1:::sub::D;GSTM1:::sub::D;NQO1:::sub::D|S22A2:::sub::D;COPT1:::sub::D;S22A3:::sub::D;ABCG2:::sub::D;MRP2:::sub::D;ATP7B:::sub::D;ATP7A:::sub::D|
Cinchocaine|ok_vet|LMNA::::8.15:C;SCN1A::::5.85:C;CP1A2::::5.3:C;CP2D6::::5.1:C;AL1A1::::5.05:C;CALM1:::inh::D;SCN5A:::inh::D;SCNAA:::inh::D|CHLE:::inh::D||
Lercanidipine|ok_inv|CCG1:::inh::D|CP2D6:::inh::D;CP3A5:::sub::D;CP3A4:::inh::D;CP3A7:::sub::D||
Foscarnet|ok|DPOL::HCMVA:inh:5.6:DC;DPOL::HHV11:inh::D||MOT1:::sub::D;S22A6:::inh::D|
Erlotinib|ok_inv|ERBB2::::10.:C;EGFR:::ant:10.:DC;ERBB2:L858R:::9.52:C;EGFR:G719S::ant:9.28:DC;EGFR:G719C::ant:9.07:DC;EGFR:L858R::ant:9.01:DC;EGFR:L861Q::ant:8.92:DC;GAK::::8.51:C;STK10::::7.72:C;M3K19::::7.6:C;SLK::::7.59:C;VGFR2::::7.3:C;ABL1:H396P:::7.24:C;ABL1:T315I:::7.23:C;ABL1:Q252H:::7.21:C;ABL1:E255K:::7.2:C;ABL1:M351T:::7.18:C;ABL1:Y253F:::7.12:C;ABL1::::7.12:C;MP2K5::::7.02:C;FLT3:D835Y:::6.89:C;EGFR:T790M::ant:6.85:DC;ABL1:F317L:::6.82:C;LYN::::6.8:C;BLK::::6.72:C;EGFR:L858R-T790M::ant:6.72:DC;ABL2::::6.7:C;ERBB4::::6.64:C;TBA1A::RAT::6.64:C;LCK::::6.6:C;FRK::::6.5:C;RET:M918T:::6.48:C;FLT3:D835H:::6.46:C;RIPK2::::6.39:C;EPHA6::::6.36:C;KC1E::::6.3:C;FLT3:N841I:::6.3:C;TNI3K::::6.24:C;AURKC::::6.22:C;TNK1::::6.2:C;ULK3::MOUSE::6.2:C;CTRO::::6.17:C;MKNK1::::6.16:C;JAK3::::6.15:C;SRC::::6.15:C;EPHA5::::6.15:C;VGFR3::::6.1:C;DDR1::::6.1:C;AURKB::::6.1:C;FLT3::::6.09:C;TIE1::::6.07:C;LTK::::6.05:C;ULK3::::6.04:C;EPHA8::::6.03:C;HIPK4::::6.02:C;MYLK2::::6.01:C;MERTK::::6.01:C;MET::::6.:C;MKNK2::::6.:C;PI42C::::6.:C;MET:Y1235D:::5.96:C;ERBB3::::5.96:C;EPHB1::::5.96:C;ABL1:F317I:::5.96:C;FGR::::5.96:C;AAK1::::5.92:C;SBK1::::5.92:C;ALK::::5.92:C;BMP2K::::5.92:C;KIT:V559D-T670I:::5.89:C;MINK1::::5.89:C;E2AK2::::5.89:C;DYRK2::::5.89:C;FLT3:K663Q:::5.89:C;RET::::5.89:C;EPHA7::::5.85:C;PGFRB::::5.85:C;KIT:D816V:::5.8:C;VGFR1::::5.8:C;KSYK::::5.8:C;KIT::::5.77:C;EPHB6::::5.77:C;HCK::::5.74:C;PGFRA::::5.74:C;FGFR2::::5.72:C;COQ8A::::5.72:C;PLK4::::5.72:C;MK09::::5.7:C;AURKA::::5.66:C;EPHB4::::5.66:C;YES::::5.66:C;M3K3::::5.64:C;EPHA3::::5.62:C;TYK2::::5.62:C;KPCD2::::5.6:C;MK04::::5.6:C;COQ8B::::5.6:C;M3K2::::5.6:C;PKN2::::5.6:C;SIK2::::5.59:C;MET:M1250T:::5.55:C;DMPK::::5.54:C;LRRK2::::5.54:C;KIT:V559D:::5.51:C;TBK1::::5.51:C;MRCKG::::5.47:C;KC1D::::5.46:C;KIT:L576P:::5.46:C;TTK::::5.43:C;JAK2::::5.43:C;TXK::::5.42:C;TYRO3::::5.41:C;UFO::::5.4:C;MK10::::5.37:C;E2AK4::::5.36:C;STK36::::5.36:C;TNIK::::5.35:C;LRRK2:G2019S:::5.32:C;RIPK4::::5.31:C;DAPK3::::5.22:C;ST17A::::5.2:C;KCC2D::::5.19:C;KS6A4::::5.15:C;GRK4::::5.14:C;SRPK3::::5.08:C;ST17B::::5.03:C;CSK::::5.02:C;LMNA::::5.:C;MRP2::::5.:C;NR1I2:::ago::D|CP3A4:::inh:5.2:DC;UD11:::inh::D;CP1B1:::sub::D;CP2C8:::inh::D;CP2D6:::sub::D;CP1A1:::sub::D;CP1A2:::sub::D;CP3A5:::sub::D|SO2B1:::inh:6.28:DC;MDR1:::sub::D;ABCG2:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Cyclophosphamide|ok_inv|NPSR1::::5.4:C;NR1I2;DNA:::cov::D|CP3A5:::sub::D;CP2C8:::sub_ind::D;CP2CI:::sub::D;CP2A6:::sub::D;CP2CJ:::sub::D;CP2B6:::sub_ind::D;CP3A4:::sub_ind::D;CP2C9:::sub::D||
Mephenytoin|ok_out|NR1I2:::act::D;SCN5A:::inh::D|CP2C9:::sub::D;CP2C8:::sub::D;CP2D6:::sub::D;CP1A2:::sub::D;CP2B6:::sub::D;CP2CJ:::inh::D||THBG:::sub::D
Rofecoxib|ok_out|PGH2:::inh:9.:DC;PGH2::MOUSE::7.92:C;PGH2::SHEEP::6.52:C;PGH2::BOVIN::6.37:C;PGH2::RAT::6.12:C;AL1A1::::5.55:C;IMPA1::RAT::5.05:C;ELN|PGH1:::sub:5.77:DC;CP2C9:::sub::D;CP2C8:::inh::D;CP3A4:::sub_ind::D;CP1A2:::inh::D|MRP4:::inh::D|
Chlormerodrin|ok_out|S12A1:::ind::D;SSDH:::inh::D|||
Cefdinir|ok|CTDS1::::5.35:C;Peptidoglycan_transpeptidase::UNK:inh::D;PERM:::inh::D;PBP3::HAEIF:inh::D;PBP2::NEIGO:inh::D||S22A8:::sub::D;S22A6:::sub::D;S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|
Guanidine|ok|ARGI::BACCD:::D;ALDH2;ENLYS::BPT4:::D;DLG4;DNA;RNAS1;GAMT;ASSY::ECOLI:::D||S47A2;S47A1:::sub::D;S22A4:::inh::D;S22A8:::inh::D;S22A5:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|
Ciprofloxacin|ok_inv|HRH3::RAT::9.18:C;TOP2A:::inh:7.52:DC;GYRB::ECOLI::6.82:C;GBRP::RAT::6.39:C;PARC::STAAU::6.:DC;LMNA::::5.25:C;AL1A1::::5.:C;GYRA::STAAU:::D;Gyrase_A::MYCTX:::D;Multidrug_resistance_protein_MdtK::ECOLX:::D;GYRA::BACSU:::D;PARE::BACSU:::D;GYRA::ECOLI:::D;KCNH2;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D;CP1A2:::inh::D|S47A2:::inh::D;S47A1:::inh::D;MDR1:::sub::D|ALBU:::bin::D
Gadoversetamide|ok_inv||||
Toremifene|ok_inv|5HT6R::::5.38:C;SHBG;ESR1:::mod::D|CP1A1:::sub::D;CP3A4:::inh::D|MDR1:::sub::D|
Nortriptyline|ok|ADA1A::RAT::10.4:C;HRH1::RAT::10.3:C;SC6A2:::inh:8.5:DC;HRH1:::ant:8.23:DC;SC6A4:::inh:8.16:DC;5HT2C:::ant:8.09:DC;ACM4:::ant:7.89:DC;5HT2A:::ant:7.82:DC;ACM5:::ant:7.7:DC;ACM1:::ant:7.7:DC;ADA2C::::7.52:C;LMNA::::7.45:C;ACM3:::ant:7.44:DC;ADA2B::::7.37:C;DRD3::::7.21:C;5HT2B::::7.07:C;ADA1B::RAT::6.94:C;ACM2:::ant:6.91:DC;ADA1D:::ant:6.87:DC;ACM1::RAT::6.8:C;5HT3A::RAT::6.77:C;5HT6R:::bin:6.67:DC;DRD1::::6.57:C;ADA2A,ADA2B,ADA2C:::ant:6.56,7.37,7.52:DC;ADA2A::::6.56:C;5HT1A::RAT::5.97:C;SC6A3::::5.88:C;5HT1B::RAT::5.84:C;RET::::5.82:C;CP2DQ::RAT::5.72:C;HRH2::::5.64:C;HRH2::CAVPO::5.15:C;TSHR::::5.1:C;5HT2C::RAT:ant::D;PGRC1,SGMR1:::bin::D;DRD2:::ant::D;ADRB1,ADRB2,ADRB3:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;5HT1A:::ant::D|CP2CJ:::sub:6.5:DC;CP2D6:::inh:6.:DC;CP1A2:::sub:5.1:DC;CP2E1:::inh::D;PGH1:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D||A1AG1;ALBU
Vincristine|ok_inv|LMNA::::8.96:C;HD::::7.75:C;TBA1A::PIG::6.66:C;TBB4B::::6.3:C;TBB2B::BOVIN::5.74:C;TBA4A:::inh::D;TBB5:::inh::D|CP3A4:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|SO1B3:::inh:5.01:DC;SO1B1:::inh::D;RBP1:::sub::D;ABCG2:::sub::D;ABCBB:::sub::D;MRP2:::inh::D;MRP7:::inh::D;MRP1:::inh::D;S22A3:::inh::D;MRP3:::inh::D;MDR1:::duo::D|
Benazepril|ok_inv|ACE:::inh:8.77:DC;ACE::RAT::8.77:C;ACE::RABIT::8.7:C|MTHR:::sub::D|S15A2:::sub::D;S15A1:::sub::D|
Amoxapine|ok|5HT2A:::ant:9.35:DC;5HT2C:::ant:8.7:DC;LMNA::::8.3:C;5HT2B:::ant:8.18:DC;TYDP1::::8.:C;HRH1:::ant:7.96:DC;SC6A2:::inh:7.89:DC;SC6A4:::inh:7.74:DC;DRD4:::ant:7.47:DC;5HT6R:::ant:7.46:DC;DRD3:::ant:7.34:DC;ADA1B::RAT::7.22:C;DRD2:::ant:7.17:DC;ADA1A::RAT::6.84:C;ADA1D::::6.82:C;DRD1:::ant:6.71:DC;5HT1A:::ant:6.66:DC;ACM4::::6.62:C;ADA2B::::6.59:C;ACM1,ACM2,ACM3,ACM4,ACM5:::ant:6.54,6.03,6.42,6.62,6.21:DC;ACM1:::ant:6.54:DC;ACM3::::6.42:C;ADA2C::::6.34:C;ADA2A,ADA2B,ADA2C:::ant:6.31,6.59,6.34:DC;ADA2A:::ant:6.31:DC;5HT7R:::ant:6.3:DC;ACM5::::6.21:C;ACM2::::6.03:C;ACM1::RAT::5.4:C;CP1A2::::5.4:C;HIF1A::::5.1:C;SMN::::5.05:C;CP3A4::::5.:C;TPO::::5.:C;SC6A3:::bin::D;GABAR:::bin::D;HRH4:::bin::D;5HT1B:::ant::D;5HT3A:::ant::D;ADA1A,ADA1B,ADA1D:::ant:,,6.82:DC;GBRA1:::ant::D;ADA1A:::ant::D|CP2D6:::inh:5.4:DC||A1AG1
Fluorouracil|ok|LMNA::::7.95:C;TPO::::7.9:C;TYSY::MOUSE::7.7:C;TSHR::::6.1:C;HD::::5.7:C;PMP22::::5.32:C;TAU::::5.25:C;END4::ECOLI::5.05:C;RNA:::destbz::D;DNA:::destbz::D|PUR1:::sub::D;UMPS:::sub::D;MTHR:::sub::D;CP2C8:::sub::D;CP2A6:::sub::D;UPP2:::sub::D;UPP1:::sub::D;DPYD:::sub::D;TYPH:::sub::D;CP1A2:::sub::D;CP2C9:::inh::D;TYSY:::sub::DC|MRP5:::sub::D;MRP4:::sub::D;MRP3:::sub::D;ABCG2:::sub::D;S29A1:::sub::D;S22A7:::sub::D|THBG:::ind::D;ALBU
Pyridostigmine|ok_inv|ACES::BOVIN::7.3:C;ACM1::RAT::7.2:C;ACES::TETCF::7.09:C;CHLE:::ant:5.46:DC;ALBU;ACES:::ant::D|||
Adinazolam|exp|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA5:::pot::D;GBRG1:::pot::D;GBRG2:::pot::D;GBRG3:::pot::D;GBRB1:::pot::D;GBRB2:::pot::D;GBRB3:::pot::D;GBRD:::pot::D;GBRE:::pot::D;GBRP:::pot::D;GBRR1:::pot::D;GBRR2:::pot::D;GBRR3:::pot::D|CP2CJ:::sub::D;CP3A4:::sub::D||
Desoximetasone|ok|GCR:::ago:8.93:DC;LMNA::::8.6:C;HIF1A::::8.3:C;NR1I2::RAT::5.:C|||
Azelaic_acid|ok|NFKB1::::8.55:C;LMNA::::8.3:C;FFP::BACIU::5.5:C;TSHR::::5.2:C;DPO1::ECOLI:inh::D;TYRO:::inh::D;S5A2:::inh::D;AK1D1:::inh::D;TRXB::STAAM:inh::D|||
Zafirlukast|ok_inv|CLTR1::CAVPO::9.52:C;CLTR1:::ant:9.52:DC;MK14::::6.45:C;MK01::::6.27:C;NR1I2::::6.15:C;AA3R::::6.11:C;S47A1::::5.89:C;STRP::STRP1::5.69:C;THAS::::5.42:C;MK03::::5.36:C;EGFR::::5.24:C;CLTR2::::5.13:C;S47A2::::5.12:C;S22A2::::5.01:C;NPSR1::::5.:C|CP2C9:::inh:5.65:DC;CP2E1:::inh::D;CP2CJ:::inh::D;CP1A2:::inh::D;CP3A4:::inh::D;PGH1:::sub::D;CP2C8:::inh::D|ABCG2:::ant::D|
Propylthiouracil|ok_inv|PERT:::inh:5.47:DC;TSHR::::5.:C|PERM:::inh:5.55:DC;CP1A1:::ind::D;DOPO:::inh::D||
Acetohydroxamic_acid|ok|MMP12:::inh::D;URE1::KLEAE:inh::D|||
Pentostatin|ok_inv|ADA::BOVIN::11.:C;ADA:::inh:10.48:DC|||
Methoxsalen|ok|ACES::::6.12:C;CP2CJ::::5.3:C;CP2D6::::5.3:C;MK01::::5.3:C;CP3A4::::5.2:C;DNA:::itc::D|CP1A2:::inh:7.8:DC;CP2AD:::inh:7.4:DC;CP2A6:::inh:6.6:DC;CP1A1:::inh::D||
Piroxicam|ok_inv|BLM::::8.05:C;NFKB1::::8.:C;PGH2::RAT::7.:C;CP3A4::::5.9:C;PGH1:::inh:5.89:DC;ACM1::RAT::5.5:C;CP2CJ::::5.2:C;PGH2:::inh::D|CP2C9:::sub:5.4:DC;CP2C8:::sub::D|S22A8:::inh:5.31:DC;SO2B1:::inh::D;S22AB:::inh::D;S22A6:::inh::D|ALBU
Lamotrigine|ok_inv|ACM1::RAT::5.6:C;CP2D6::::5.2:C;SCN2A:::inh:5.:DC;5HT3A:::inh::D;5HT2A:::inh::D;ACM1,ACM2,ACM3,ACM4,ACM5:::inh::D;OPRK:::inh::D;HRH1:::inh::D;GBRA1,GBRA2,GBRA3,GBRA4,GBRA5,GBRA6,GBRG1,GBRG2,GBRG3:::inh::D;GABAR:::inh::D;DRD2:::inh::D;DRD1,DRD5:::inh::D;ADRB1:::inh::D;ADA2A:::inh::D;ADA1A:::inh::D;AA2AR:::inh::D;AA1R:::inh::D;CAC1E:::inh::D|UD11:::sub_ind::D;UD13:::sub::D;DYR:::inh::D;UD14:::sub::D|S22A2:::inh::D;MDR1:::sub::D|
Perflutren|ok||||
Hydroxyzine|ok|HRH1:::ant::D|CP3A5:::sub::D;CP3A4:::sub::D;CP2D6:::inh::D||
Zanamivir|ok_inv|NRAM::INBLE::10.:C;NRAM::I34A1::9.3:C;NRAM::I33A0::9.1:C;NRAM::I68A0::8.58:C;NEUR2:::inh:5.28:DC;NEUR3::::5.17:C;NRAM::INBBE:inh::D;NRAM::I79A0:inh::D|||
Bosentan|ok_inv|EDNRA::RAT::8.33:C;EDNRA:::ant:8.33:DC;EDNRA::PIG::8.12:C;EDNRB:::ant:7.1:DC;EDNRB::RAT::7.02:C;NR1I2::::5.05:C|CP2C9:::sub_ind::D;CP3A4:::sub_ind::D|ABCBB:::inh::D|
Tigecycline|ok|RS19::ECOLI:cov::D;RS14::ECOLI:cov::D;RS13::ECOLI:cov::D;RS12::ECOLI:cov::D;RS9::ECOLI:cov::D;16S_ribosomal_RNA::Gut_flora:cov::D|||
Doxapram|ok_vet|CP2D6::::7.:C;KCNK9:::inh::D;KCNK3:::inh::D|||
Benzthiazide|ok|CP2C9::::5.4:C;CAH12:::inh::D;CAH9:::inh::D;CAH4:::inh::D;CAH2:::inh::D;CAH1:::inh::D;S12A3:::inh::D|||
Methotrexate|ok|DYR::RAT::10.14:C;DRTS::LEIMA::9.89:C;DYR::PNECA::9.:C;DYR::STAAU::9.:C;DYR::LACCA::8.89:C;DYR::ENTFC::8.85:C;DRTS::TOXGO::8.85:C;DYR::BOVIN::8.77:C;LMNA::::8.35:C;DYR::MOUSE::8.18:C;DYR::MYCTU::8.08:C;DYR::CHICK::7.72:C;PTR1::LEIMA::7.41:C;P53::::7.:C;NCOA3::::6.68:C;TYSY::LACCA::5.3:C;TAU::::5.:C;LOX15::::5.:C|DYR:::sub:10.42:DC;TYSY:::sub:6.22:DC;FOLC:::sub:5.49:DC;CP3A4:::sub::D;GGH:::sub::D;6PGD:::inh::D;MTHR:::sub::D;AOXA:::sub::D;PUR9:::inh::DC|S19A1:::sub:7.92:DC;FOLR2:::sub:6.97:DC;FOLR1:::sub:6.94:DC;PCFT:::inh:6.92:DC;S36A1:::sub::D;S15A1:::sub::D;SO4C1;SO1B1:::sub::D;S22A7:::sub::D;ABCG2:::sub::D;SO3A1:::sub::D;SO1C1:::sub::D;S22AB:::sub::D;SO1B3:::sub::D;ABCCB:::sub::D;MOT1:::sub::D;SO1A2:::sub::D;MDR1:::sub::D;MRP2:::inh::D;S22A8:::inh::D;MRP7:::inh::D;S22A6:::inh::D;MRP1:::inh::D;MRP4:::inh::D;MRP3:::inh::D|ALBU:::bin::D
Carbamazepine|ok_inv|LMNA::::8.4:C;TSHR::::5.2:C;NR1I2:::act::D;ACHA4;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A:::inh::D|UD17:::ind::D;UD16:::ind::D;UD11:::ind::D;UD2B7:::sub::D;CP3A5:::sub_ind::D;CP2B6:::sub_ind::D;CP2CJ:::duo::D;CP2C9:::ind::D;CP1A2:::duo::D;CP2C8:::sub_ind::D;CP3A4:::sub_ind::D|MRP2:::sub::D;RBP1:::sub::D;MDR1:::ind::D|
Cisatracurium|ok|LMNA::::6.9:C;CP3A4::::5.:C;ACHA2:::ant::D|||
Succimer|ok|Lead:::chel::D;Mercury:::chel::D;Cadmium:::chel::D;Arsenic:::chel::D|||
Cephalexin|ok_inv_vet|MK01::::5.1:C;PBPA::STRR6:inh::D;PBP2::STRR6:inh::D;PBP1B::STRR6:inh::D;PBP2A::STRR6:inh::D;PBP3::STREE:inh::D||S22A8:::inh::D;S47A1:::sub::D;S22A6:::inh::D;S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|ALBU
Cinnarizine|ok_inv|LMNA::::8.3:C;HRH1:::ant:8.06:DC;SGMR1::::7.77:C;DRD3::::7.07:C;ADA2C::::7.02:C;5HT2A::::6.99:C;ACM3::::6.79:C;ADA2A::::6.78:C;DRD2::::6.59:DC;SCN1A::::6.36:C;5HT2B::::6.33:C;ADA1B::RAT::6.3:C;ACM4::::6.29:C;ACM5::::6.26:C;ADA1D::::6.24:C;SC6A4::::6.24:C;ACM1,ACM2,ACM3,ACM4,ACM5:::bin:6.22,,6.79,6.29,6.26:DC;ACM1::::6.22:C;5HT1A::RAT::6.21:C;ADA1A::RAT::6.11:C;OPRM::::6.04:C;ADA2B::::5.99:C;SC6A3::::5.88:C;ACM1::RAT::5.75:C;END4::ECOLI::5.75:C;SC6A2::::5.55:C;DRD1,DRD5:::bin::D;CAC1I:::inh::D;CAC1H:::inh::D;CAC1G:::inh::D;CAC1S:::inh::D;CAC1F:::inh::D;CAC1D:::inh::D;CAC1C:::inh::D|CP3A4:::sub:5.5:DC;CP1A1:::sub::D;CP2A6:::sub::D;CP2B6:::sub::D;CP1A2:::sub::D;CP2C9:::sub::D;CP2D6:::sub::D||
Fondaparinux|ok_inv|FA10:::inh::D;ANT3:::pot::D|||
Vinblastine|ok|TBB4B::::7.15:C;TBB::PIG::6.22:C;TBB2B::BOVIN::6.22:C;THAS::::5.73:C;LOX15::RABIT::5.3:C;MDR1B::MOUSE::5.1:C;JUN;TBE:::cov::D;TBG1:::cov::D;TBD:::cov::D;TBB5:::cov::D;TBA1A:::cov::D|CP2D6:::inh::D;CP3A4:::duo::D|MDR1:::duo:7.:DC;SO1B1:::inh::D;ABCBB:::inh::D;MRP6:::inh::D;MRP2:::duo::D;MRP1:::duo::D|
Propranolol|ok_inv|ADRB2:::ant:9.62:DC;ADRB2::CAVPO::9.01:C;ADRB1:::ant:8.9:DC;ADRB2::CANLF::8.75:C;ADRB1::RAT::8.62:C;ADRB1:W134A:RAT::8.:C;ADRB1:Y356F:RAT::7.5:C;ADRB1:S190A:RAT::7.4:C;5HT1B::RAT::7.3:C;5HT1A::RAT::7.05:C;ADRB3:::ant:7.:DC;ADRB1:Y356A:RAT::6.7:C;SC6A4::::6.69:C;5HT2B::::6.66:C;5HT2A::::6.38:C;5HT2C::::5.92:C;SGMR1::::5.92:C;5HT6R::::5.85:C;SCN5A::::5.68:C;KCNH2::::5.55:C;5HT1A::::5.4:DC;NTCP::::5.26:C;5HT1B|CP2D6:::inh:5.72:DC;CP1A2:::sub:5.4:DC;AOFA:::inh::D;CP1A1:::inh::D;CP3A4:::sub::D;CP2CJ:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|MDR1:::sub::D;S22A2:::inh::D|ALBU;A1AG1
Atropine|ok_vet|ACM4:::ant:9.98:DC;ACM3::RAT::9.92:C;ACM5:::ant:9.68:DC;ACM1:::ant:9.6:DC;ACM1::RAT::9.59:C;ACM3:::ant:9.49:DC;ACM2:::ant:9.46:DC;ACES::MOUSE::9.46:C;ACM2::MOUSE::9.46:C;ACM4::RAT::9.28:C;ACM2::RAT::9.15:C;ACM5::RAT::9.07:C;5HT2C::::6.28:C;ADA1D::::6.18:C;ACHB2;ACHA4;GLRA1:::ant::D||ABCBB:::sub::D|
Fenoprofen|ok|PGH1:::inh:6.84:DC;PPARG;PPARA:::act::D;PGH2:::inh::D|||ALBU
Fenfluramine|ok_ill_inv_out|TAU::::6.9:C;5HT2A;5HT2C:::ago::D;5HT2B:::ago::D;SC6A4:::inh::D|CP2D6:::inh::D||
Clonidine|ok|ADA2A::RAT::9.41:C;ADA2C::RAT::8.82:C;ADA2A::BOVIN::8.7:C;ADA2A:::ago:8.42:DC;ADA2B:::ago:8.21:DC;ADA2B::RAT::8.08:C;NISCH::::8.05:C;ADA2C:::ago:8.03:DC;NISCH::RAT::7.85:C;ADA1A::BOVIN::7.05:C;ADA1B::RAT::6.94:C;ADA1A::RAT::6.82:C;LMNA::::6.55:C;ADA1A:::ago:6.54:DC;S22A1::::6.26:C;ADA1D:::ago:6.23:DC;S22A1::RAT::5.85:C;5HT1A::RAT::5.51:C;5HT1A::::5.49:C;CP2CJ::::5.3:C;CP2C9::::5.1:C;ADA1B:::ago::D|CP2D6:::sub:5.1:DC;CP3A5:::sub::D;CP1A1:::sub::D;CP3A4:::sub::D;CP1A2:::sub::D|MDR1:::sub::D;S22A4:::inh::D;S22A5:::inh::D;S22A3:::inh::D|ALBU:::bin::D
Sulfamethizole|ok_inv_vet|LMNA::::5.35:C;DHPS::ECOLI:inh::D|CP2C9:::inh::D||ALBU
Valaciclovir|ok_inv|AMPC::ECOLI::5.55:C;KITH::HHV1:sub::D;DPOL::HHV11:inh::D|KITH::HHV1C:sub::D;KGUA:::sub::D|NTCP2:::sub::D;S6A14;S22A6;S22A8:::sub::D;S15A2:::inh::D;S15A1:::inh::D|
Carbenicillin|ok_inv|DACA,DACB,DACC,PBPA,PBPB,MRDA,FTSI::ECOLI:inh::D|PA24A:::inh::D|S22A6:::inh::D|
Mazindol|ok_inv|SC6A2:::inh:8.31:DC;SC6A3::RAT::8.15:C;SC6A3:::inh:7.66:DC;SC6A4:::inh:7.3:DC;SC6A4::RAT::6.64:C;SGMR1::::6.63:C;VMAT2|||
Valdecoxib|ok_out|PGH2:::inh:8.3:DC;CAH12::::7.89:C;CAH9::::7.57:C;CAH2:::inh:7.37:DC;CAN::CANAL::7.37:C;CAH15::MOUSE::7.18:C;CAH5B::::7.06:C;CAH14::::6.97:C;CAH::METTE::6.89:C;CAH4::BOVIN::6.47:C;CAH13::MOUSE::6.37:C;CAH13::::6.37:C;CAH6::::6.24:C;CAN::YEAST::6.18:C;MTCA2::MYCTU::6.17:C;CAH5A::::6.04:C;COX2::::5.96:C;CAH4::::5.87:C;SC6A2::::5.54:C;CAH7::::5.41:C;CAH3:::inh::D|UD19:::sub::D;CP2C9:::inh::D;CP3A4:::sub::D||
Lactulose|ok|BGA2::ECOLI:::D|||
Voriconazole|ok|CP51::CANAL:ant::D|CP2B6:::inh:6.47:DC;CP2C9:::inh:5.55:DC;CP2CJ:::inh:5.29:DC;PGH1:::sub::D;CP3A4:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;FMO3:::sub::D;FMO1:::sub::D||
Levocarnitine|ok_inv|AMPC::ECOLI::5.85:C;PERM;EST1;XDH;CPT1A:::act::D;CPT2;OCTC;MCAT;MCATL;CACP||S22A8:::sub::D;S22AG:::sub::D;SO1B1:::inh::D;S22A5:::sub::DC;S22A4:::inh::DC|
Enalapril|ok_vet|ACE:::inh:8.92:DC;ACE::RABIT::8.7:C;LMNA::::7.65:C;ACE::RAT::6.85:C||SO1A2:::sub::D;S22A7:::inh::D;S22A8:::inh::D;S22A6:::inh::D;S15A1:::inh::D;MDR1:::inh::D|ALBU:::bin::D
Nizatidine|ok|HRH2:::ant::D|CHLE:::inh::D|MDR1:::sub::D|
Diclofenac|ok_vet|PGH1:::inh:8.52:DC;PGH1::BOVIN::8.52:C;PGH2:::inh:8.3:DC;IL8::::8.1:C;CXCR1::::7.92:C;PGH2::MOUSE::7.66:C;PGH2::SHEEP::7.22:C;PGH1::SHEEP::7.17:C;PGH2::RAT::6.3:C;AK1BA::::5.72:C;FABPL::RAT::5.49:C|PA2GA:::inh::D;LOX5:::pot::D;UD2B4:::sub::D;UD19:::sub::D;UD13:::sub::D;CP2E1:::inh::D;CP2CI:::sub::D;CP2B6:::sub::D;CP3A4:::inh::D;UD2B7:::sub::D;CP2C8:::sub::D;CP1A2:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D|S22A6:::inh:5.4:DC;KCNQ3:::ago::D;KCNQ2:::ago::D;ASIC1:::inh::D;SCN4A:::inh::D;ABCBB:::sub::D;SO1B1:::inh::D;SO1C1:::inh::D;S22AB:::inh::D;S22A8:::inh::D;MRP1:::inh::D;MRP4:::inh::D|TTHY::::6.:DC;ALBU::::5.61:DC
Fluticasone_propionate|ok|GCR:::ago:10.12:DC;GCR::RAT::9.12:C;MCR:::ant::D;PA24A:::inh::D;PRGR:::ago::D|CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::inh::D;CP3A4:::inh::D||SO1B1:::inh::D;MDR1:::sub::D;CBG
Lisuride|ok_inv|DRD3:::ago:10.23:DC;ADA2A::::9.94:DC;ADA2B::::9.63:DC;5HT1A::RAT::9.58:C;DRD2:S194A:RAT::9.52:C;DRD2:S197A:RAT::9.4:C;5HT1A:::ago:9.4:DC;DRD2:::ago:9.3:DC;DRD2::RAT::9.22:C;ADA2C::::9.2:DC;5HT2A:::ago:9.06:DC;5HT2B:::ant:8.49:DC;5HT1B::RAT::8.34:C;5HT6R::::8.26:C;ADA1A::RAT::8.04:C;5HT2C:::ago:8.:DC;CP2D6::::7.8:C;HRH1::::7.72:C;ADA1D::::7.7:C;ADRB2::::7.54:C;ADA1B::RAT::7.17:C;DRD1:::ant:7.11:DC;ADRB1::::6.49:C;HRH2::::5.99:C;5HT7R;5HT1B:::ago::D;5HT1D:::ago::D;DRD5:::ant::D;DRD4:::ago::D|CP3A4:::sub::D||
Doxazosin|ok|ADA1B::RAT::9.51:C;ADA1A:::ant:9.27:DC;ADA1A::RAT::9.2:C;ADA1B::::9.13:DC;ADA1D:::ant:9.09:DC;ADA1D::RAT::8.97:C;5HT4R::CAVPO::6.9:C;SC6A3::::6.83:C;5HT2B::::6.63:C;5HT2C::::6.55:C;ADA2C::::6.55:C;KCNH2,KCNH6,KCNH7:::inh:6.23,,:DC;KCNH2::::6.23:C;ADA2A::::6.14:C;SC6A4::::5.85:C;ADRB2::::5.72:C;MMP1::::5.24:C|CP2C9:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D;CP2CJ:::sub::D|S22A1:::inh::D;MDR1:::inh::D|
Fluocinolone_acetonide|ok_inv_vet|HIF1A::::8.89:C;GCR:::ago:8.85:DC;MK01::::5.5:C;ANXA5:::ind::D;ANXA4:::ind::D;ANXA3:::ind::D;ANXA2:::ind::D;ANXA1:::ind::D|CP3A4:::sub_ind::D||CBG:::bin::D
Piperazine|ok_vet|GBRB3:::ago::D|CP2D6:::sub::D||
Ethosuximide|ok|RORG::MOUSE::5.55:C;CAC1G:::inh::D|CP3A4,CP343,CP3A5,CP3A7:::sub::D;CP3A4:::sub::D;CP2E1:::sub::D||
Amiloride|ok|LMNA::::6.15:C;SCNNA:::inh:6.11:DC;SL9A2::RABIT::6.:C;SL9A1::RAT::6.:C;UROK:::inh:5.6:DC;AA2AR:H250N:::5.48:C;AOFA::::5.41:C;ASIC3::::5.36:C;S22A2::RAT::5.33:C;HCD2::::5.3:C;S22A1::RAT::5.16:C;AOC3::RAT::5.:C;SL9A1:::inh::D;ASIC1:::inh::D;ASIC2:::inh::D;SCNND:::inh::D;SCNNG:::inh::D;SCNNB:::inh::D|AOC1::PIG:inh::D;AOC1:::inh::DC|S22A4:::inh::D;S22A2:::inh::D|
Oxytetracycline|ok_inv_vet|TYDP1::::6.4:C;DPOLB::::5.55:C;MEN1::::5.45:C;TAU::::5.2:C;HIF1A::::5.1:C;16S_ribosomal_RNA::Gut_flora:inh::D;RS4::ECOLI:inh::D;RS9::ECOLI:inh::D||S22A7:::inh::D;S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D|
Ulobetasol|ok|GCR:::ago::D|||CBG
Gadoteridol|ok_inv||||
Labetalol|ok|ADRB1:::ant:8.23:DC;ADRB2:::ant:7.96:DC;ADA1A::RAT::7.64:C;ADRB2::CAVPO::7.4:C;ADA1A,ADA1B,ADA1D:::ant:6.8,,6.59:DC;ADA1A::::6.8:C;5HT1A::RAT::6.65:C;ADA1D::::6.59:C;ADA1B::RAT::6.49:C;SGMR1::::6.12:C;SC6A3::::5.89:C;5HT2B::::5.71:C;SC6A2::::5.48:C|CP2D6:::inh:6.1:DC;UD19:::sub::D;UD2B7:::sub::D;UD11:::sub::D;CP2CJ:::sub::D|ABCB5|A1AG1,A1AG2:::sub::D;ALBU:::sub::D
Thiopental|ok_vet|CAC1C::CAVPO::6.55:C;LMNA::::6.45:C;ACM3;FAAH1:::inh::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2CJ:::sub::D;CP3A4,CP343,CP3A5,CP3A7:::sub::D||
Monobenzone|ok|PGH1::::5.99:C;CP1A2::::5.8:C;PGH2::::5.43:C;SC6A2::::5.41:C;LOX15::RABIT::5.31:C;CP2CJ::::5.2:C;HIF1A::::5.:C;FRIL::HORSE::5.:C;LMNA::::5.:C;TYRO:::inh::D|||
Linezolid|ok_inv|STRP::STRP1::6.8:C;23S_ribosomal_RNA::Gut_flora:inh::D|AOFB:::inh:5.68:DC;AOFA:::inh:5.1:DC||
Ivermectin|ok_inv_vet|GLRA2::RAT::6.67:C;NR1H4::::6.59:C;AA3R::::6.54:C;MDR1B::MOUSE::6.3:C;MDR1A::MOUSE::6.3:C;ADA2C::::6.24:C;DRD3::::6.12:C;ACM1::::5.92:C;ACM3::::5.89:C;ADA2A::::5.66:C;DRD1::::5.65:C;ACM5::::5.59:C;SC6A3::::5.45:C;SC6A2::::5.41:C;AT1A2::RAT::5.19:C;AT2A2::RAT::5.17:C;AT1A1::RAT::5.08:C;GBRB3:::ago::D;GLRA3:::ago::D|CP3A4:::sub_ind::D|MDR1:::inh:7.97:DC;MRP1:::inh:6.3:DC;SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::sub::D;MRP2:::inh::D|
Medroxyprogesterone_acetate|ok_inv|PRGR:::ago:10.:DC;ANDR::::8.54:C;ANDR::RAT::8.32:C;ANDR::MOUSE::8.21:C;GCR::::8.06:C;AK1C3::::6.55:C;SHBG::::6.2:C;AK1C1::::6.15:C;ESR2::::6.03:C;MCR::::5.92:C;AK1C2::::5.8:C;NPSR1::::5.6:C;GABAR:::inh::D;MDR1:::inh::D;ESR1:::ago::D|CP3A1::RAT:sub::D;CP2C9:::inh::D;3BHS2:::inh::D;CP2C8:::inh::D;CP3A4:::sub_ind::D||ALBU:::bin::D
Cisapride|ok_out|5HT4R:::ago::D;5HT3A:::ago::D;5HT2A:::ago::D;KCNH2:::inh::D|CP3A7:::sub::D;CP3A4:::sub::D;CP3A5:::sub::D;CP2A6:::sub::D;CP2B6:::sub::D;CP2CJ:::inh::D;CP2C8:::sub::D;CP2C9:::inh::D;CP2D6:::inh::D||
Sulindac|ok_inv|LMNA::::8.25:C;MK01::::7.4:C;CP2CJ::::6.7:C;ALDR:::inh:6.43:DC;GLRA1::::6.42:C;ALDR::RAT::6.36:C;CP3A4::::6.2:C;CP1A2::::5.4:C;PGH2:::inh:5.06:DC;AK1BA:::inh::D;PD2R2:::ant::D;PPARD:::neg::D;MK03:::inh::D;PGH1:::inh::D|CP1A1:::inh::D|S22A6:::inh::D|ALBU
Cyclothiazide|ok|THB::::6.85:C;GRIA1::::6.:C;GRIA2::::5.65:C;GRIA4::::5.42:C;GRIA2::RAT::5.21:C;LMNA::::5.2:C;SFRP4:::inh::D;CAH4:::inh::D;CAH2:::inh::D;CAH1:::inh::D;ATNG:::inh::D||S22A6:::inh::D|
Nafcillin|ok_inv|PBPA::STRR6:inh::D;PBP3::STREE:inh::D;PBP2A::STRR6:inh::D;PBP2::STRR6:inh::D;PBP1B::STRR6:inh::D|CP1A2:::ind::D;CP3A4:::ind::D|S22A6:::inh::D|ALBU
Chloroquine|ok_inv_vet|HRP1::PLAFA::7.12:C;NQO2::::5.82:C;RBP::CHICK::5.68:C;KCNH2::::5.6:C;PRIO::::5.4:C;GST::PLAFA:inh::D;TLR9;TNFA;Fe_II_protoporphyrin_IX::PLAFA:ant::D;GSTA2|CP3A5:::sub::D;CP2C8:::sub::D;CP1A1:::sub::D;CP2D6:::inh::D;CP3A4:::sub::D|MDR1:::inh::D|
Ethionamide|ok|PPO2::AGABI::5.4:C;KATG::MYCTU:::D;INHA::MYCTU:cov::D|||
Metaraminol|ok_inv|ADA1A:::ago::D|||
Butorphanol|ok_ill_vet|OPRK:::ago:9.92:DC;OPRM:::antp:9.92:DC;OPRD:::ago:7.92:DC|||
Bisoprolol|ok|ADRB2:::ant::D;ADRB1:::ant::D|CP3A4:::sub::D|MDR1:::inh::D|
Amodiaquine|ok_inv|CP2J2::::6.:C;HNMT:::inh::D;Fe_II_protoporphyrin_IX::PLAFA:cov::D|CP2D6:::inh:6.19:DC;CP2C9:::inh::D;CP1B1:::sub::D;CP1A1:::sub::D;CP2C8:::sub::D|MDR1:::inh::D|
Furazolidone|exp_vet|RORG::MOUSE::6.3:C;P53::::5.:C;DNA:::cov::D|AOFA:::inh::D;AOFB:::inh::D||
Rifabutin|ok_inv|ENPL;HS90A;RPOC::ECOLI:inh::D;RPOB::ECOLI:inh::D;RPOA::ECOLI:inh::D|CP2C9:::ind::D;CP2C8:::ind::D;CP2B6:::ind::D;CP2CJ:::ind::D;CP3A4:::sub_ind::D|MDR1:::ind::D|
Paramethadione|ok|CAC1I:::sup::D|CP2E1:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D||
Demeclocycline|ok|RS4::ECOLI:inh::D;RS9::ECOLI:inh::D|||
Imatinib|ok|DDR1:::ant:9.15:DC;ABL1:::inh:8.96:DC;ABL1:Q252H::inh:8.74:DC;PGFRA:::ant:8.7:DC;ABL1:F317L::inh:8.6:DC;ABL1:H396P::inh:8.23:DC;ABL2::::8.22:C;ABL1:F317I::inh:8.08:DC;ABL1:M351T::inh:8.07:DC;ABL1::MOUSE::7.97:C;CSF1R:::ant:7.96:DC;KIT:::ant:7.89:DC;KIT:L576P::ant:7.85:DC;PGFRB:::ant:7.85:DC;KIT:V559D::ant:7.82:DC;DDR2::::7.82:C;KIT:A829P::ant:7.82:DC;CAH2::::7.52:C;CAH1::::7.5:C;NQO2::::7.41:C;LCK::::7.4:C;S47A1::::7.4:C;ABL1:Y253F::inh:7.36:DC;KIT:V559D-V654A::ant:7.15:DC;CAH9::::7.12:C;ABL1:E255K::inh:7.11:DC;CAH15::MOUSE::7.11:C;KIT:K642E::ant:7.01:DC;CAH7::::6.96:C;PGFRB::RAT::6.79:C;THAS::::6.7:C;LYN::::6.7:C;PGFRB::MOUSE::6.52:C;FRK::::6.5:C;ABL1:T315I::inh:6.47:DC;S47A2::::6.46:C;ABL1:G250E::inh:6.44:DC;PI42C::::6.42:C;CAH6::::6.41:C;CAH14::::6.33:C;CAH3::::6.28:C;BLK::::6.28:C;5HT2A::::6.27:C;KIT:D816H::ant:6.25:DC;SC6A4::::6.13:C;KIT:D816V::ant:6.09:DC;HIPK4::::6.02:C;CAH12::::6.01:C;MK10::::6.:C;GAK::::6.:C;IRAK1::::5.92:C;CLK4::::5.9:C;EPHA8::::5.85:C;RAF1::::5.77:C;MELK::::5.72:C;HRH2::::5.71:C;FGR::::5.62:C;CYSP::TRYCR::5.6:C;KIT:V559D-T670I::ant:5.6:DC;M3K20::::5.59:C;SRC::CHICK::5.56:C;ST17A::::5.55:C;FYN::::5.51:C;MK08::::5.49:C;BRAF:V600E:::5.48:C;TAOK1::::5.4:C;TNI3K::::5.37:C;CLK1::::5.35:C;CAH4::::5.34:C;KSYK::::5.3:C;MK09::::5.28:C;CDK19::::5.26:C;FLT3::::5.2:C;CAH13::MOUSE::5.13:C;EGFR::::5.12:C;PLK4::::5.11:C;TYK2::::5.06:C;NTRK1:::ant::D;RET_proto_oncogene:::inh::D;BCR:::inh::D|CP2C8:::sub::D;PGH1:::sub::D;CP2CJ:::sub::D;CP2D6:::inh::D;CP2C9:::inh::D;CP1A2:::sub::D;CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D|ABCG2:::inh:6.3:DC;S22A2:::inh:5.38:DC;MDR1:::inh:5.14:DC;ABCBB:::sub::D;ABCA3:::sub::D;S22A1:::sub::D|A1AG1:::sub::D;ALBU:::sub::D
Triamcinolone|ok_vet|BLM::::8.35:C;LMNA::::7.65:C;GCR:::ago:7.59:DC;NFKB1::::7.55:C;HIF1A::::7.5:C;CP2J2::::5.02:C|CP3A7:::sub_ind::D;CP3A5:::sub_ind::D;CHLE:::ind::D;PGH2:::inh::D;CP3A4:::sub_ind::D||ALBU:::bin::D;CBG:::bin::D
Oxandrolone|ok_inv|ANDR:::ago::D|CP2C9:::inh::D||
Nicardipine|ok_inv|CAC1C::RAT::9.08:C;CAC1C:::inh:6.6:DC;TRPA1::MOUSE::6.3:C;ADA2C::RAT::5.85:C;CP2J2::::5.77:C;LMNA::::5.7:C;MDR1A::MOUSE::5.6:C;AA3R::::5.49:C;ADA1B::RAT::5.44:C;S29A1::RAT::5.27:C;MDR1B::MOUSE::5.1:C;TAU::::5.05:C;CALM1;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;ADA1D:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;PDE1B:::inh::D;PDE1A:::inh::D;CAC1D:::inh::D;CA2D1:::inh::D;CACB2:::inh::D|CP2C9:::inh:6.55:DC;CP3A4:::inh:6.42:DC;CP2CJ:::inh:6.25:DC;CP2C8:::inh:5.81:DC;CP2D6:::inh:5.8:DC;CP3A5:::inh::D;CP2E1:::sub::D;CP2B6:::ind::D|MDR1:::inh:6.02:DC;ABCBB:::sub::D;SO1B1:::inh::D|
Fluphenazine|ok|DRD3::::9.69:C;DRD2:::ant:9.27:DC;5HT2A::::8.84:DC;HRH1::::8.33:C;SGMR1::::8.07:C;ADA1A::RAT::8.02:C;DRD1:::ant:7.96:DC;ADA2B::::7.89:C;ADA1D::::7.8:C;ADA1B::RAT::7.72:C;DRD5::::7.68:C;ADA2C::::7.66:C;5HT6R::::7.62:C;5HT2B::::7.6:C;5HT2C::::7.46:DC;ADA2A::::7.1:C;ACM4::::6.32:C;ACM1::::6.19:C;ANDR::RAT::6.1:C;SC6A4::::6.1:C;5HT1B::RAT::6.06:C;5HT1A::RAT::6.03:C;ACM3::::6.:C;CP1A2::::6.:C;HRH2::::5.92:C;SC6A3::::5.79:C;PDR5::YEAST::5.77:C;SC6A2::::5.71:C;DRD4::::5.69:C;ACM2::::5.58:C;LMNA::::5.45:C;SCN1A::::5.43:C;KCNH2::::5.33:C;KCNK2::::5.33:C;AA3R::::5.17:C;ACM1::RAT::5.15:C;NK2R::::5.13:C;FYN::::5.1:C;OPRM::::5.07:C;OPRD::::5.07:C;MC5R::::5.05:C;OPRK::::5.:C;ANDR;CALM1:::inh::D|CP2D6:::inh:6.2:DC;CP2E1:::inh::D|MDR1:::inh:5.24:DC|
Testosterone|ok_inv|ANDR::RAT::8.85:C;ANDR::MOUSE::8.7:C;ANDR:::ago:8.57:DC;TSHR::::7.5:C;CAC1C::::7.47:C;CBG::::6.72:C;SGMR1::::5.92:C;GCR::::5.84:C;S5A1::RAT::5.72:C;SO1A1::RAT::5.27:C;LMNA::::5.25:C;ERG2::YEAST::5.11:C;MCR:::lig::D;ESR1:::inh::D|CP19A:::sub:6.22:DC;CP3A4:::sub_ind:5.:DC;CP2C8:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP2B6:::sub::D;CP2AD:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D;CP11A:::inh::D;AOFA:::ind::D;CP343:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|SO1B3:::sub::D;ABCG2:::sub::D;NTCP:::inh::D;S22A7:::inh::D;S22A8:::ind::D|SHBG:::bin:9.2:DC;ALBU:::bin::D
Efavirenz|ok_inv|NPSR1::::5.:C;Reverse_transcriptase_RNaseH::9HIV1:inh::D|UD11:::ind::D;CP2C8:::inh::D;CP2D6:::inh::D;CP1A2:::inh::D;CP3A7:::ind::D;CP3A5:::ind::D;CP3A4:::duo::D;CP2B6:::duo::D;CP2C9:::inh::D;CP2CJ:::duo::D|S22A1:::inh::D;ABCBB:::sub::D|ALBU
Bacitracin|ok_vet|5HT1B::RAT::5.87:C;LCK::::5.72:C;EGFR::::5.27:C;A2MG:::inh::D;IDE:::inh::D;C55_isoprenyl_pyrophosphate::G+-Bac:ant::D||BCRC::BACLI:sub::D;BCRB::BACLI:sub::D;BCRA::BACLI:sub::D|
Niacin|ok_inv_nutra|HCAR2:::ago:8.06:DC;AA3R::::8.:C;HCAR2::MOUSE::7.54:C;HCAR2::RAT::7.48:C;LYAG::::5.45:C;S6A11::RAT::5.22:C;SC6A1::MOUSE::5.1:C;SC6A1::::5.1:C;NNMT:::bin::D;NADC:::bin::D;HCAR3:::ago::D|CP2E1:::inh::D;CP3A4:::inh::D;CP2D6:::inh::D|MOT4;SC5A8;MOT1:::sub::D;SO2B1:::inh::D;S22A5:::inh::D|THBG:::inh::D
Clorazepic_acid|ok_ill|TSPO:::ago::D;GABAR:::aga::D|CP3A4:::sub::D||
Guanabenz|ok_inv|ADA2C::RAT::8.77:C;ADA2A:::ago:7.82:DC;NISCH::::7.46:C;5HT2B::::7.21:C;ADA2B:::bin:7.17:DC;TAAR1::::7.05:C;5HT2C::::6.97:C;5HT2A::::6.95:C;ADA1A::RAT::6.8:C;ADA2C::::6.79:C;ADA1D::::6.63:C;ADA1B::RAT::6.35:C;5HT1A::RAT::5.93:C;AOFA::::5.75:C;MTOR::::5.68:C|CP1A2:::sub::D||
Alendronic_acid|ok|FPPS:::inh:7.35:DC;VATA:::inh::D;PTPRE:::inh::D;PTPRS:::inh::D;PTN4:::inh::D;Hydroxylapatite:::ant::D|||
Clofarabine|ok_inv|DNA;RIR1:::inh::D;DPOLA:::inh::D|DCK:::sub::D|ABCG2:::sub::D|
Docosanol|ok_inv|VGP3::EBVP3:itc::D;GP350::EBVB9:itc::D|||
Dexmedetomidine|ok_vet|ADA1D::::10.82:C;ADA2C::RAT::10.82:C;ADA2A::RAT::10.82:C;ADA2C::::9.32:C;ADA2A:::ago:9.1:DC;ADA1B::RAT::8.3:C;CP3A4::::6.8:C;CP2C9::::6.7:C;ADA1A::BOVIN::6.42:C;CP2CJ::::5.3:C|CP1A2:::inh:6.8:DC;CP2D6:::inh::D;CP1A1:::inh::D;CP2E1:::sub::D||
Sulfacetamide|ok|TSHR::::6.2:C;FOL1::YEAST:inh::D;DHP1::ECOLX:inh::D;DHPS::ECOLI:inh::D|||
Prednisone|ok_vet|GCR:::ago:6.28:DC;RORG::MOUSE::5.45:C;AL1A1::::5.:C|DHI1:::sub::D;CP2C9:::ind::D;CP2C8:::ind::D;CP2B6:::ind::D;CP1B1:::ind::D;CP2A6:::ind::D;CP3A4,CP343,CP3A5,CP3A7:::ind::D;CP3A5:::ind::D;CP2CJ:::ind::D;CP3A4:::sub_ind::D|SO1A2:::inh::D;MDR1:::sub_ind::D|CBG:::bin::D;ALBU:::sub::D
Clofibrate|ok_inv|ACM1::RAT::8.2:C;TSHR::::5.6:C;AMPC::ECOLI::5.25:C;FABPL::RAT::5.22:C;PPARA:::ago::D|CP3A4:::sub_ind:5.:DC;CP4AB:::sub_ind::D;CP1A1:::ind::D;GSTA2:::inh::D;CP2E1:::ind::D||THBG:::ind::D
Astemizole|ok_out|KCNH2:::inh:9.05:DC;HRH1:::ant:8.79:DC;FNTA::BOVIN::8.7:C;HRH1::CAVPO::8.42:C;5HT2A::::8.25:C;5HT2B::::8.13:C;ADA1A::RAT::8.:C;5HT2C::::7.03:C;ADA1B::RAT::7.02:C;DRD3::::6.83:C;ACM3::::6.75:C;ACM1::::6.59:C;ACM4::::6.59:C;ADA2C::::6.55:C;ADA1D::::6.42:C;5HT1A::RAT::6.36:C;ACM2::::6.3:C;ACM5::::6.3:C;OPRM::::6.22:C;5HT1B::RAT::6.2:C;SC6A4::::6.15:C;SC6A3::::6.1:C;SGMR1::::6.03:C;NK2R::::6.:C;CAC1C::::5.96:C;MDR1A::MOUSE::5.89:C;SC6A2::::5.87:C;DRD2::::5.82:C;5HT6R::::5.82:C;TAU::::5.8:DC;HRH2::::5.78:C;MDR1B::MOUSE::5.77:C;ADA2B::::5.76:C;ADA2A::::5.74:C;DRD1::::5.7:C;DRD4::::5.67:C;MC5R::::5.67:C;RORG::MOUSE::5.6:C;OPRK::::5.58:C;FYN::::5.55:C;MEN1::::5.5:C;SSR5::::5.39:C;GLRA1::::5.38:C;OPRD::::5.34:C;ADRB3::::5.22:C;EGFR::::5.22:C;CP2CJ::::5.1:C;HRH4::::5.1:C;LMNA::::5.1:C;CP1A2::::5.1:C;NK1R::::5.06:C;ADRB1::::5.:C;KCNH1|CP3A4:::inh:5.48:DC;CP2D6:::sub:5.1:DC;CP2J2:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|MDR1:::inh:6.52:DC;ABCBB:::sub::D|
Inulin|ok_inv_nutra|Cycloinulo_oligosaccharide_fructanotransferase::PAEMA:bin::D|||
Butoconazole|ok|Ergosterol::CANAL:::D|||
Adenosine|ok_inv|AA3R:::ago:8.94:DC;AA1R:::ago:8.63:DC;AA2BR::RAT::8.3:C;AA1R::RAT::8.29:C;AA2AR:::ago:7.7:DC;AA2AR::RAT::7.52:C;AA2BR:::ago:7.29:DC;AA3R::RAT::7.:C;STAT6::::5.9:C;S28A1::::5.74:C;AA1R::CAVPO::5.47:C;S28A2::::5.28:C;ADK::TOXGO::5.05:C|ADK:::sub::D;ADA:::sub::D|S28A3::::5.68:DC|
Simvastatin|ok|HMDH:::inh:8.59:DC;HMDH::RAT::8.37:C;CHLE::HORSE::6.12:C;ACES::ELEEL::5.74:C;HDAC2:::inh::D;ITAL:::inh_allo::D|CP2C8:::inh:5.43:DC;CP2CJ:::sub::D;UD2B7:::sub::D;UD13:::sub::D;UD11:::sub::D;CP2B6:::duo::D;CP2D6:::sub::D;CP2C9:::inh::D;CP3A5:::sub::D;CP3A4:::sub::D|SO1B1:::inh:5.36:DC;MDR1:::inh:5.05:DC;SO1B3;SO2B1;ABCBB:::sub::D;MRP2:::sub::D;SO1A2:::inh::D|
Pemetrexed|ok_inv|TYSY:::inh:8.89:DC;DYR:::inh:8.15:DC;PUR2:::inh:7.93:DC;PCFT::::7.88:C;FOLR1::::7.38:C;FOLR2::::7.22:C;S19A1::::6.86:C;TYSY::MOUSE::6.47:C;DRTS::TOXGO::6.37:C;TYSY::LACCA::6.26:C;DYR::MOUSE::6.25:C;DYR::LACCA::5.64:C;PUR9:::inh::D|S29A1:::ind::D;DCK:::ind::D|S22A8:::sub::D|
Mebendazole|ok_vet|HIF1A::::6.1:C;LMNA::::6.05:C;LEF::BACAN::5.6:C;VGFR2::::5.44:C;CP1A2::::5.4:C;ABL1::::5.34:C;HD::::5.25:C;TBB4B:::inh::D;TBA1A:::inh::D|CP3A4,CP343,CP3A5,CP3A7:::sub::D;CP1A1:::ind::D||
Gonadorelin|ok_inv_vet|GNRR2:::ago::D;GNRHR:::ago::D|||
Dyclonine|ok|IMPA1::RAT::8.89:C;AL1A1::::6.65:C;LMNA::::6.2:C;CP2C9::::5.6:C;CP1A2::::5.5:C;CP2D6::::5.3:C;LEF::BACAN::5.3:C;RORG::MOUSE::5.:C;SCNAA:::inh::D|||
Nystatin|ok_vet|Ergosterol::CANAL:bin::D||SO1B3:::inh::D;SO1B1:::inh::D|
Dextropropoxyphene|ok_ill_inv_out|EST1;OPRK:::ant::D;OPRD:::ago::D;OPRM:::ago::D|CP2D6:::inh::D;CP3A4:::inh::D||
Mitotane|ok|BLM::::7.65:C;5HT6R::::6.19:C;SC6A3::::6.1:C;SC6A2::::6.09:C;SC6A4::::5.8:C;ADA2A::::5.56:C;5HT2B::::5.51:C;AA3R::::5.38:C;TAU::::5.3:C;LMNA::::5.2:C;ANDR:::ant::D;PRGR;ESR1;ADX;C11B1:::ind::D|CP3A4:::ind::D||THBG:::ind::D;CBG;SHBG
Stavudine|ok_inv|BLM::::6.1:C;ACM1::RAT::5.55:C;Reverse_transcriptase_RNaseH::9HIV1:inh::D||S28A1;S22A6:::sub::D|ALBU
Leucovorin|ok|DYR::::5.63:C;SO1A3::RAT::5.09:C||S22A8:::inh::D|
Dyphylline|ok|PDE7B:::inh::D;PDE7A:::inh::D;AA2AR:::ant::D;AA1R:::ant::D;PDE4D:::inh::D;PDE4C:::inh::D;PDE4A:::inh::D;PDE4B:::inh::D|||
Pentazocine|ok_vet|SGMR1::CAVPO::8.66:C;SGMR1:::ago:8.51:DC;OPRM::RAT::8.16:C;SGMR1::RAT::7.92:C;OPRK::CAVPO::7.12:C;OPRK:::ago::D;OPRM:::ant::D|||
Magnesium_sulfate|ok_inv_vet|CCG1;CA2D1;CAC1C;CACB1;CACB2;CAC1S|||
Latanoprost|ok_inv|TAU::::5.3:C;PF2R:::ago::D|Corneal_esterases:::sub::D|S22A8:::inh::D;S22A6:::inh::D;SO2A1:::sub::D|
Estrone|ok|ESR1:::ago:9.15:DC;HCD2::::8.89:C;ESR2::::8.68:DC;DHB1::::8.52:C;SHBG::::8.18:DC;LMNA::::7.95:C;HIF1A::::7.8:C;BLM::::6.7:C;CP19A::::5.6:DC;PMP22::::5.57:C;SC6A4::::5.55:C;NFKB1::::5.4:C;LOX15::RABIT::5.18:C;ANDR::RAT::5.11:C;5HT2B::::5.06:C;CBG::::5.:C;ANDR|CP1A2:::sub:5.9:DC;CP3A4:::sub:5.7:DC;CP3A5:::sub::D;CP2E1:::sub::D;CP2C9:::sub::D;CP2B6:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D|ABCG2:::inh:5.52:DC;S22A8:::sub::D;SO1B1:::inh::D;SO1A2:::inh::D;MDR1:::sub_ind::D;SO2B1:::inh::D|ALBU
Trazodone|ok_inv|5HT2A:::ant:8.25:DC;5HT2A::RAT::7.77:C;HRH1:::ant:7.38:DC;5HT2C:::ago:7.33:DC;ADA1A::RAT::7.33:C;ADA1B::RAT::7.21:C;5HT2B::::7.17:C;SC6A4:::inh:6.99:DC;ADA1D::::6.89:C;5HT1A::RAT::6.75:C;ADA2B::::6.75:C;ADA2C::::6.55:C;ADA2A:::ant:6.47:DC;5HT1B::RAT::6.08:C;SGMR1::::6.03:C;DRD3::::5.9:C;ALBU::RAT::5.1:C;5HT2C::RAT:ant_pago::D;ADA1A:::ant::D;5HT1A:::ant_pago::D|CP2D6:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|MDR1:::ind::D|
Mecamylamine|ok_inv|ACHB2;ACHA4;ACHA7;ACHA2:::ant::D|||
Sevelamer|ok|Phosphate:::bin::D|||
Acamprosate|ok_inv|GRM5:::ant::D;NMDA:::ant::D;GABAR:::ago::D||S36A1|
Metaxalone|ok||||
Verapamil|ok|CAC1C::RAT::8.85:C;TSPO::RAT::8.85:C;KCNH2:::inh:8.:DC;CAC1S::RAT::7.24:C;DRD3::::7.2:C;CAC1C::CAVPO::7.:C;5HT2B::::6.98:C;5HT2A::::6.9:C;SC6A4::::6.9:DC;CAC1C:::inh:6.82:DC;5HT2C::::6.81:C;ADA2A::::6.66:C;ADA1A::RAT::6.07:C;ADA1B::RAT::6.03:C;ADA1A:::ant:6.:DC;CAC1C::RABIT::6.:C;5HT1A::RAT::5.76:C;MDR1B::MOUSE::5.7:C;HRH2::::5.59:C;SCN1A::::5.48:C;KCNA3::::5.1:C;MDR1A::MOUSE::5.:C;ADA1D:::ant::D;ADA1B:::ant::D;CAC1H:::inh::D;CAC1G:::inh::D;KCJ11:::inh::D;CAC1A:::inh::D;CAC1B:::inh::D|CP3A4:::inh:5.33:DC;CP2D6:::inh::D;CP2E1:::sub::D;CP1A2:::sub::D;CP2CJ:::sub::D;CP2B6:::act::D;CP2CI:::sub::D;CP3A5:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D|MDR1:::inh:7.54:DC;S22A1:::inh:5.54:DC;MRP1:::inh:5.46:DC;S47A2:::inh::D;S47A1:::inh::D;MRP7:::inh::D;MRP4:::inh::D;SO1A2:::inh::D;SO1B1:::inh::D;MRP3:::inh::D;S22A5:::inh::D;S22A4:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Trimethobenzamide|ok_inv|LMNA::::7.25:C|||
Flumethasone|ok_vet|HIF1A::::8.3:C;RAB9A::::6.:C;RORG::MOUSE::5.05:C;GCR:::ago::D|CP3A4:::sub::D||CBG:::bin::D
Sulfametopyrazine|ok_out|Dihydropteroate_synthetase::PLAFA:inh::D|||
Nilutamide|ok_inv|ACM1::RAT::8.8:C;ANDR:::ant:8.05:DC;TSHR::::6.9:C;LMNA::::5.75:C;CP1A2::::5.6:C;CP3A4::::5.4:C;LOX12::::5.2:C;NFKB1::::5.15:C;RORG::MOUSE::5.05:C|CP2CJ:::inh:6.9:DC;NCPR:::sub::D||
Nafarelin|ok|GNRR2:::ago::D;GNRHR:::ago::D|||
Epinephrine|ok_vet|ADA2A:::ago:8.3:DC;ADA2C::RAT::7.89:C;ADRB2::CAVPO::7.82:C;ADA1B::RAT::7.77:C;ADRB3::::7.51:C;ADRB2:::ago:6.71:DC;ADA1D:::ant:6.66:DC;ADRB1::RAT::6.64:C;ADA1A::RAT::6.6:C;ADA2C::::6.45:C;ADA2B:::ago:6.4:DC;ADA1A:::ago:6.4:DC;ADRB2::CANLF::6.18:C;ADRB2::RAT::6.14:C;HCD2::::6.1:C;DRD2::::6.04:C;HIF1A::::5.8:C;TYDP1::::5.5:C;LOX15::RABIT::5.48:C;OPRM::RAT::5.4:C;MK01::::5.4:C;KDM4E::::5.15:C;FFP::BACIU::5.15:C;TAU::::5.1:C;TNFA:::duo::D;ADRB1:::ago::D;ADA1B:::ago::D|AOFA,AOFB:::sub::D;COMT:::sub::D;CP3A4:::inh::D;CP2C9:::inh::D|S22A1:::sub::D;S22A2:::sub::D|
Sumatriptan|ok_inv|5HT1B:::ago:9.3:DC;5HT1D:::ago:8.92:DC;5HT1B::GORGO::8.19:C;5HT2C::::8.14:C;5HT1B::RAT::8.09:C;5HT3A::::8.03:C;5HT1D::PIG::7.7:C;5HT1F:::ago:7.59:DC;5HT1D::RAT::7.21:C;5HT1A:::ago:6.64:DC;5HT2A::::6.42:C;5HT1A::MOUSE::6.35:C;5HT1A::RAT::6.34:C;5HT5A::::6.3:C;5HT1E::::5.26:C;S47A1::::5.17:C|AOFA:::sub::D|SO1B1:::sub::D;ABCG2:::sub::D;MDR1:::sub::D;SO1A2:::ind::D|
Pirenzepine|ok|ACM4::::8.94:C;ACM1:::ant:8.83:DC;ACM1::RAT::8.42:C;AA3R::::7.66:C;ACM3::RAT::7.55:C;ACM4::RAT::7.46:C;ACM5::::7.45:C;ACM3::::7.32:C;ACM2::RAT::6.92:C;LMNA::::6.9:C;ACM2::::6.76:C;ACM1::DROME::6.41:C;ACM5::MOUSE::6.12:C;CP1A2::::5.1:C|||
Cefixime|ok_inv|PLCG1::::5.92:C;APAF::::5.04:C;MRDA::HAEIN:inh::D||S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|
Chlorpropamide|ok_inv|LMNA::::8.3:C;NFKB1::::6.35:C;TSHR::::5.8:C;THB::::5.7:C;NPSR1::::5.3:C;ABCC8:::inh::D|PGH1:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D|S22A6:::inh::D;S15A2:::inh::D;S15A1:::inh::D|
Aprepitant|ok_inv|NK1R:::ant:10.1:DC;NK1R::MERUN::10.05:C;NK3R::::6.34:C|CP3A4:::duo:7.34:DC;CP2C9:::duo::D;CP2CJ:::inh::D||
Galantamine|ok|ACES:::inh:7.21:DC;CHLE:::inh:6.77:DC;ACES::ELEEL::6.44:C;ACES::TETCF::6.44:C;ACES::RAT::6.27:C;ACES::MOUSE::5.68:C;CHLE::HORSE::5.49:C;ACES::BOVIN::5.06:C;ACHB4:::alo::D;ACHB3:::alo::D;ACHB2:::alo::D;ACH10:::alo::D;ACHA9:::alo::D;ACHA7:::alo::D;ACHA6:::alo::D;ACHA5:::alo::D;ACHA4:::alo::D;ACHA3:::alo::D;ACHA2:::alo::D;ACHE:::alo::D;ACHG:::alo::D;ACHD:::alo::D;ACHB:::alo::D;ACHA:::alo::D|CP2D6:::sub::D;CP3A4:::sub::D||
Tamoxifen|ok|ESR2:::duo:9.29:DC;EBP:::inh:9.:DC;EBPL::::8.55:C;ESR1:::duo:8.1:DC;SGMR1::::8.06:C;PRGR::::6.89:C;ERR1::::6.7:C;5HT2C::::6.62:C;DRD3::::6.44:C;ACM3::::6.2:C;ACM1::::6.17:C;ACM4::::6.17:C;ADA2A::::6.14:C;KCNH2:::inh:6.1:DC;THAS::::6.04:C;5HT6R::::5.98:C;FYN::::5.92:C;NK2R::::5.91:C;SC6A4::::5.91:C;5HT2B::::5.88:C;5HT2A::::5.86:C;SC6A2::::5.84:C;SC6A3::::5.84:C;ERG2::YEAST::5.82:C;ADA2B::::5.79:C;ACM5::::5.73:C;AA3R::::5.68:C;ADA1D::::5.61:C;ACM2::::5.56:C;ERBB2::::5.53:C;EGFR::::5.45:C;DRD4::::5.41:C;AA2AR::::5.4:C;DRD1::::5.37:C;PGH1::::5.36:C;OPRD::::5.33:C;DRD2::::5.33:C;AMPC::ECOLI::5.3:C;ADRB3::::5.24:C;STRP::STRP1::5.21:C;OPRK::::5.2:C;5HT1A::RAT::5.16:C;OPRM::::5.15:C;LCK::::5.1:C;NK1R::::5.07:C;ADA1A::RAT::5.05:C;HRH2::::5.03:C;ADRB1::::5.:C;MK08:::mod::D;SHBG:::ind::D;ERR3;NR1I2;ANDR;KPCA,KPCB,KPCD,KPCE,KPCG,KPCI,KPCT,KPCZ:::inh::D|CP3A4:::duo:6.7:DC;CP2B6:::inh:6.05:DC;ST1E1:::sub::D;UDB17:::sub::D;UD2B7:::sub::D;CP1A2:::sub::D;ST2A1:::sub::D;ST1A1:::sub::D;UD110:::sub::D;CP2E1:::sub::D;CP2A6:::sub::D;CP19A:::inh::D;EST1:::inh::D;CP2C8:::inh::D;FMO3:::sub::D;FMO1:::sub::D;CP1B1:::inh::D;CP1A1:::sub::D;CP2CJ:::sub::D;CP2C9:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP2D6:::inh::D|MDR1:::duo:7.:DC;ABCA1:::sub::D;ABCBB:::inh::D;MRP2:::sub::D;ABCG2:::sub::D|THBG:::ind::D;ALBU:::sub::D
Benzyl_benzoate|ok|LIPS::RAT::5.96:C|||
Isoflurophate|ok_out|EST1::PIG::7.3:C;ACES:::inh:6.92:DC;ACES::ELEEL::6.32:C;PPGB::::5.:C;TRFE|CHLE:::inh::DC||ALBU
Losartan|ok|AGTR1:::ant:9.48:DC;AGTR1::RABIT::8.8:C;AGTRB::RAT::8.74:C;AGTRA::RAT::8.17:C;AGTR1::CAVPO::7.74:C;ACE::::7.72:C;AGTR2::::7.72:C;AGTR1::BOVIN::7.02:C;SO1B1::::6.8:C;SO1B3::::6.05:C;AGTR2::RAT::5.13:C|CP2C9:::sub:5.54:DC;CP2C8:::inh::D;UDB17:::sub::D;UD2B7:::sub::D;UD110:::sub::D;UD13:::sub::D;UD11:::sub::D;CP2CJ:::inh::D;CP3A4:::inh::D|ABCBB:::sub::D;GTR9:::inh::D;S22AC:::inh::D;S22A6:::inh::D;MDR1:::inh::D|ALBU:::sub::D
Thioridazine|ok_out|5HT2A:::ant:8.9:DC;ACM1::::8.77:C;ACM1::RAT::8.7:C;ADA1A::RAT::8.69:C;ADA1B::RAT::8.59:C;DRD2::RAT::8.55:C;ADA1D::::8.54:C;DRD3::::8.47:C;ACM5::::8.18:C;HRH1::::8.08:C;ACM4::::7.96:C;DRD2:::ant:7.92:DC;DRD1::RAT::7.76:C;5HT2B::RAT::7.74:C;ACM3::::7.72:C;5HT2C::::7.64:C;ADA2C::::7.6:C;KCNH2:::inh:7.48:DC;5HT6R::::7.48:C;5HT1A::RAT::7.47:C;ACM2::::7.42:C;ADA2A::::7.3:C;5HT7R::::7.15:C;5HT2B::::7.09:C;DRD5::RAT::7.07:C;DRD1:::ant:7.01:DC;HRH1::RAT::7.:C;SGMR1::::6.82:C;ADA2B::::6.76:C;SC6A4::::6.4:C;DRD4::::6.29:C;SGMR1::RAT::6.12:C;HRH2::::6.03:C;OPRK::::6.:C;PDR5::YEAST::5.89:C;CAC1C::CAVPO::5.89:C;ADA2C::RAT::5.89:C;CAC1C::::5.88:C;SC6A2::::5.81:C;SCN5A::::5.74:C;SC6A3::::5.72:C;EGFR::::5.53:C;FYN::::5.3:C;SCN1A::::5.19:C;ALBU::RAT::5.17:C;PIM1::::5.16:C;5HT1B::RAT::5.06:C;CP1A2::::5.03:C;ADA1B:::ant::D;ADA1A:::ant::D|CP2D6:::inh:5.75:DC;CP2CJ:::sub:5.2:DC;CP2E1:::inh::D||
Moricizine|ok_out|HIF1A::::5.8:C;CP3A4::::5.3:C;SCN5A:::inh::D|||
Amphotericin_B|ok_inv|LMNA::::7.1:C;CYSP::TRYCR::5.1:C;Ergosterol::CANAL:bin::D|CP3A4:::inh::D||
Warfarin|ok|AMPC::ECOLI::5.45:C;ALBU::RAT::5.03:C;NR1I2;VKOR1:::inh::D|CP2CI:::sub::D;CP2C8:::inh::D;CP3A4:::sub_ind::D;CP2CJ:::inh::D;CP1A2:::sub::D;CP2C9:::sub_ind::D||ALBU::::5.7:DC;A1AG1
Midazolam|ok_ill|GBRP::RAT::8.7:C;TSPO::RAT::8.7:C;S22A1::::5.43:C;GBRA6:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA5:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP3A4:::inh:5.61:DC;CP3A7:::sub::D;UD14:::sub::D;CP3A5:::sub::D||
Tobramycin|ok_inv|16S_ribosomal_RNA::Gut_flora:inh::D;RS12::ECOLI:inh::D|AAC2::MYCTU:sub::D||
Trovafloxacin|ok_out|THAS::::5.4:C;TOP2A:::inh::D;PARC::HAEIN:inh::D;GYRA::HAEIN:inh::D|CP1A2:::inh::D||
Pentosan_polysulfate|ok|FGF2:::ant::D;FGF1:::ant::D;FGF4:::inh::D|||
Fludrocortisone|ok_inv|GCR:::ago::D;MCR:::ago::D|DHI1:::sub::D;DHI2:::sub::D;CP3A4:::sub::D||CBG:::sub::D;ALBU:::sub::D
Mycophenolate_mofetil|ok_inv|PTPS:::inh::D;IMDH2:::inh::D;IMDH1:::duo::D|Q6IPK9:::sub::D;CP2C8:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D;EST1:::sub::D;UD110:::sub::D;UD18:::sub::D;UD2B7:::sub::D;UD19:::sub::D;UD16:::sub::D;UD17:::sub::D;UD11:::sub::D|MRP2;MDR1:::sub::D;ABCG2:::sub::D;SO1B3:::sub::D;SO1B1:::sub::D|
Cephaloglycin|ok|Multimodular::BACLI:ant::D||S22A5:::inh::D|
Flurazepam|ok_ill_inv|GBRT:::pot::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP3A4:::sub::D;CP2A6:::sub::D;CP2E1:::inh::D|S22A2:::inh::D;MDR1:::inh::D|
Moexipril|ok|ACE:::inh:8.59:DC;ACE2:::inh::D||S15A2:::sub::D;S15A1:::sub::D|
Phentolamine|ok|ADA1A:::ant:9.22:DC;ADA1A::BOVIN::9.1:C;ADA2A::BOVIN::9.03:C;ADA2C::RAT::8.85:C;ADA2A:::ant:8.77:DC;ADA1B::RAT::8.57:C;ADA1A::RAT::8.33:C;ADA2A::RAT::8.33:C;ADA1B:::ant:8.32:DC;ADA1A::RABIT::8.2:C;ADA1D:::ant:8.12:DC;ADA2B::::8.12:C;ADA2C::::8.08:C;NISCH::::7.94:C;ADA1D::RAT::7.35:C;5HT2A::::6.99:C;5HT2C::::6.68:C;ADA1B::MESAU::6.66:C;SGMR1::::6.26:C;CP2D6::::6.1:C;5HT2B::::5.62:C;LMNA::::5.3:C;SCN1A::::5.08:C|||
Fluorescein|ok|KV230;DNA||S22A6:::inh::D;ABCBB:::sub::D;MRP1:::sub::D|
Daunorubicin|ok|RORG::MOUSE::7.2:C;MMP2::::5.72:C;HD::::5.65:C;MEN1::::5.55:C;FFP::BACIU::5.5:C;TAU::::5.35:C;APEX1::::5.:C;TOP2B:::inh::D;TOP2A:::inh::D;DNA:::itc::D|NCPR:::sub::D;XDH:::sub::D;CP1B1:::inh::D;CP1A1:::sub::D;CP3A5:::ind::D;CP3A4:::inh::D|MRP1:::inh:7.15:DC;MDR1:::duo:5.6:DC;ABCG2:::sub::D;ABCBB:::sub::D;MRP6:::sub::D;MRP2:::inh::D;MRP7:::sub::D|
Furosemide|ok_vet|CAH14::::7.28:C;CAH1::::7.21:C;CAH2:::inh:7.19:DC;CAH6::::6.61:C;CAH12::::6.58:C;CAH5B::::6.49:C;CAH9::::6.38:C;CAH5A::::6.3:C;CAH7::::6.29:C;CAH13::MOUSE::6.26:C;CAH4::::6.25:C;CISD1::::5.64:C;GPR35:::ago:5.49:DC;DHI1::MOUSE::5.42:C;DHI1::::5.42:C;S22A6::RAT::5.02:C;S12A1:::inh::D|UD11:::sub::D;6PGD:::inh::D|S22AB:::inh::D;SO2A1:::inh::D;MRP2:::inh::D;S22A8:::inh::D;S22A5:::inh::D;S22A6:::duo::D|THBG:::bin::D;ALBU:::bin::D
Ergotamine|ok|5HT1B::RAT::10.04:C;5HT1A::RAT::9.35:C;ADA2A:::pag:9.1:DC;5HT1D:::ago:9.1:DC;5HT6R::::9.02:C;DRD2:::ago:8.84:DC;DRD3::::8.83:C;ADA2B:::ago:8.76:DC;ADA2C::::8.74:C;5HT2A:::ago:8.73:DC;5HT1B:::ago:8.68:DC;5HT2B::::8.66:DC;ADA1A::RAT::8.49:C;ADA1B::RAT::8.34:C;5HT5A::::7.85:C;ADA1D:::pag:7.62:DC;5HT2C:::ago:7.54:DC;5HT4R::CAVPO::6.58:C;DRD1,DRD5:::ago:6.06,:DC;DRD1::::6.06:C;ADRB2::::5.72:C;ADRB1::::5.62:C;THAS::::5.51:C;FYN::::5.5:C;LCK::::5.19:C;5HT1F:::ago::D;5HT1A:::ago::D;SC6A2:::inh::D;ADA1B:::pag::D;ADA1A:::pag::D|CP3A4:::inh:6.:DC|MDR1:::inh::D|
Tizanidine|ok_inv|NISCH:::ago:7.55:DC;ADA2A,ADA2B,ADA2C:::ago:7.07,,5.91:DC;ADA2A::::7.07:C;ADA1A::BOVIN::6.58:C;ADA2C::::5.91:C;ADA1A,ADA1B,ADA1D:::ago::D|CP1A2:::sub::D||
Nitrofurantoin|ok_vet|CISD1::::6.09:C;LMNA::::6.:C;LEF::BACAN::5.9:C;STRP::STRP1::5.23:C;TYDP1::::5.05:C;RS10::ECOLI:inh::D;NFSA::ECOLI:pot::D;NIFJ::ECOLI:pot::D|NCPR:::sub::D|MRP2;MDR1:::sub::D;ABCBB:::sub::D;ABCG2:::sub::D|
Nicergoline|ok_inv|ADA1A:::ant::D|CP2D6:::sub::D||
Eplerenone|ok|MCR:::ant:6.91:DC|C11B2:::inh::D;CP3A5:::sub::D;CP3A4:::sub::D||
Amprenavir|ok_inv|LMNA::::6.2:C;THAS::::5.17:C;Pol_polyprotein::9HIV1:inh::D|CP3A5:::sub:6.7:DC;CP3A4:::duo:6.59:DC;CP2D6:::sub::D;CP2C9:::sub::D;CP2CJ:::inh::D;CP2B6:::inh::D|SO1B1:::inh::D;MRP1:::inh::D;MDR1:::sub_ind::D|
Icodextrin|ok_inv||AMYP:::sub::D||
Methazolamide|ok|CAH3:::inh::D;CAH7:::inh::D;CAH2:::inh::D;CAH4:::inh::D;CAH1:::inh::D||S22A6:::inh::D|
Naltrexone|ok_inv_vet|OPRD:::ant:10.7:DC;OPRK:::ant:10.4:DC;OPRM:::ant:10.3:DC;OPRM::MOUSE::9.8:C;OPRM::CAVPO::9.77:C;OPRK::CAVPO::9.51:C;OPRM::RAT::9.34:C;SGMR1::RAT::9.3:C;OPRK::MOUSE::9.09:C;OPRK::RAT::8.97:C;OPRD::MOUSE::8.36:C;OPRD::RAT::8.32:C;CP2D6::::6.:C;HCG20471_isoform_CRA_c:::ant::D|UD11:::sub::D||
Delavirdine|ok|Reverse_transcriptase_RNaseH::9HIV1:inh::D|CP2CJ:::inh::D;CP2C9:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D||
Tamsulosin|ok_inv|ADA1D::RAT::10.6:C;ADA1A:::ant:10.54:DC;ADA1A::RAT::10.52:C;ADA1D:::ant:10.24:DC;ADA1A::BOVIN::9.9:C;ADA1B:::ant:9.89:DC;ADA1A::RABIT::9.8:C;ADA1B::MESAU::9.7:C;ADA1B::RAT::9.69:C;DRD3::::9.55:C;5HT1A::::9.1:C;ADA2B::RAT::8.17:C;ADA2C::::8.1:C;DRD2::::7.89:C;ADA2A::::7.87:C;5HT7R::::7.08:C;5HT1B::RAT::6.03:C|CP2D6:::sub::D;CP3A4:::sub::D||A1AG1
Porfimer_sodium|ok_inv|LDLR;FCGR1:::ant::D|||
Sufentanil|ok_inv|SGMR1::RAT::10.7:C;OPRM::RAT::9.66:C;MDR1::::5.35:C;OPRK;OPRD:::ago::D;OPRM:::ago::D|CP3A4:::sub::D||
Lamivudine|ok_inv|HSF1::MOUSE::6.54:C;TAU::::5.45:C;DPOL::HBVF1:inh::D;DNA:::cov::D;Reverse_transcriptase_RNaseH::9HIV1:inh::D|NT5C:::sub::D;PCY2:::sub::D;PCY1A:::sub::D;NDKB:::sub::D;NDKA:::sub::D;PGK1:::sub::D;KCY:::sub::D;DCK:::sub::D|MRP2;MRP3:::sub::D;MRP4:::sub::D;MDR1:::sub::D;S22A3:::sub::D;S22A2:::sub::D;S22A1:::sub::D;ABCG2:::sub::D;S22A6:::sub::D;MRP1:::inh::D|ALBU
Ibandronate|ok_inv|FPPS:::inh:8.44:DC;FDFT::RAT::6.19:C;Hydroxylapatite:::ant::D|||
Diethylcarbamazine|ok_inv_vet|PGH1:::inh::D;LOX5:::inh::D|CHLE:::inh::D||
Flurbiprofen|ok_inv|PGH2:::inh:8.:DC;PGH1:::inh:8.:DC;PGH1::SHEEP::7.96:C;PGH1::RAT::6.77:C;PGH2::MOUSE::6.3:C;FABPL::RAT::5.93:C;AK1C3::::5.81:C;TSHR::::5.2:C|UD2B4:::sub::D;UD19:::sub::D;UD13:::sub::D;UD11:::inh::D;UD2B7:::sub::D;CP2C9:::sub::D|S22A6:::inh:5.82:DC;MRP4:::inh::D|ALBU
Oxacillin|ok_inv|Penicillin_binding_protein_2::STAAU:::D;PBPA::CLOPE:inh::D;PBP1B::STRR6:inh::D;PBP2::STRR6:inh::D;PBPA::STRR6:inh::D;PBP2A::STRR6:inh::D;PBP3::STREE:inh::D||S15A2:::inh::DC;S15A1:::inh::DC|
Apomorphine|ok_inv|DRD2::RAT::9.4:C;DRD2:::ago:9.21:DC;DRD5::RAT::9.:C;DRD1::BOVIN::9.:C;DRD4::RAT::8.82:C;DRD1::RAT::8.77:C;DRD3:::ago:8.59:DC;DRD4:::ago:8.37:DC;DRD1:::ago:8.34:DC;HCD2::::7.7:C;DRD3::RAT::7.61:C;ADA2C::RAT::7.2:C;DRD1::MOUSE::7.:C;5HT7R::RAT::6.73:C;DRD2::BOVIN::6.7:C;TYDP1::::6.55:C;5HT1A::RAT::6.53:C;5HT1A:::ago:6.53:DC;SGMR1::RAT::6.52:C;DRD2:S197A:RAT::6.22:C;DRD2:S194A:RAT::5.92:C;PGDH::::5.4:C;5HT3A::RAT::5.35:C;CP3A4::::5.3:C;P53::::5.2:C;ADA1B::RAT::5.11:C;CP2CJ::::5.:C;CALY:::ago::D;5HT1B:::ago::D;5HT1D:::ago::D;ADA2A:::ago::D;5HT2B:::ago::D;5HT2A:::ago::D;DRD5:::ago::D;5HT2C:::ago::D;ADA2B:::ago::D;ADA2C:::ago::D|||
Paroxetine|ok_inv|SC6A4:::inh:10.4:DC;SC6A4::RAT::9.82:C;SC6A3::MOUSE::9.36:C;SC6A2::MOUSE::7.7:C;ACM4::::7.47:C;ACM1,ACM2,ACM3,ACM4,ACM5:::inh:7.46,6.72,7.42,7.47,7.05:DC;ACM1::::7.46:C;ACM3::::7.42:C;SC6A2:::inh:7.4:DC;ACM5::::7.05:C;ACM2::::6.72:C;SC6A3::::6.4:C;SC6A3::RAT::6.4:C;NK1R::::6.05:C;P2RX4::::5.73:C;SGMR1::::5.65:C;P2RX4::RAT::5.61:C;MTOR::::5.53:C;CAC1C::::5.41:C;ADA1B::RAT::5.27:C;ADA2C::RAT::5.2:C;NORA::STAAU::5.15:C;KCNH2::::5.07:C;DRD1,DRD5;5HT2B:::ago::D;5HT1A,5HT1B,5HT1D,5HT1E,5HT1F,5HT2A,5HT2B,5HT2C,5HT3A,5HT3B,5HT3C,5HT3D,5HT3E,5HT4R,5HT6R,5HT7R;HRH1:::inh::D;DRD2;ADRB1,ADRB2,ADRB3:::inh::D;ADA2A,ADA2B,ADA2C:::bin::D;ADA1A,ADA1B,ADA1D:::bin::D;5HT2A:::ago::D|CP2D6:::inh:6.:DC;CP2CJ:::inh::D;CP3A4:::inh::D;CP1A2:::inh::D;CP2B6:::inh::D;CP2C9:::inh::D|MDR1:::inh::D|
Nedocromil|ok_inv|HS90A;PD2R;FPR1:::ant::D;CLTR2:::ant::D;CLTR1:::sup::D|||
Norethisterone|ok|PRGR:::ago:9.4:DC;ESR1::RAT::9.2:C;ANDR::RAT::7.82:C;GCR:::ago:6.71:DC;ESR1::::6.64:C;SC6A4::::5.62:C;ANDR:::ago::D|CP2A6:::sub::D;CP1A2:::sub::D;CP2CJ:::sub_ind::D;AK1D1:::sub::D;S5A1,S5A2,PORED:::sub::D;3BHS2:::sub::D;AK1C4:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|SHBG:::sub:7.97:DC;ALBU:::sub::D
Adefovir_dipivoxil|ok_inv|DPOL::HBVD2:::D|NDKB:::sub::D;NDKA:::sub::D;KAD4:::sub::D;KAD2:::sub::D|S22A3:::sub::D;MRP5:::sub::D;MRP4:::sub::D;S22A6:::inh::D|
Azatadine|ok|HRH1::RAT::8.41:C;HRH1:::ant::D|CP3A4:::ind::D||
Clodronic_acid|ok_inv_vet|Hydroxylapatite:::ant::D;ADT3:::inh::D;ADT2:::inh::D;ADT1:::inh::D|PGH2:::inh::D||
Procaine|ok_inv_vet|CP2D6::::5.:C;AOFA,AOFB:::inh::D;LPP60:::inh::D;PA24A:::inh::D;KCMA1,KCMB1,KCMB2,KCMB3,KCMB4,KCNN4,KCNN1,KCNN2,KCNN3:::bin::D;DNA:::bin::D;ACHA2:::ant::D;SC6A3:::inh::D;5HT3A:::ant::D;NMD3A:::ant::D;SCNAA:::inh::D|CHLE:::inh::D||
Lisinopril|ok_inv|ACE:::inh:10.:DC;ACE::RABIT::8.22:C;RENI:::inh::D||S15A2:::sub::D;S15A1:::inh::D|
Methoxamine|ok_inv|ADA1A:::ago:6.14:DC;ADA2C::RAT::5.44:C;ADA1D:::bin::D;ADA1B:::ago::D|||
Imiquimod|ok_inv|ADA1D::::5.89:C;HRH2::::5.83:C;TLR7:::ago:5.67:DC;AA2AR::::5.52:C;TLR8:::ago::D|CP3A4:::sub::D||
Homatropine_methylbromide|ok|ACM2:::ant::D;ACM1:::ant::D;ACM4:::ant::D;ACM5:::ant::D;ACM3:::ant::D|||
Trimipramine|ok|5HT2C::RAT:bin::D;ACM1,ACM2,ACM3,ACM4,ACM5:::bin::D;ADRB1,ADRB2,ADRB3:::bin::D;DRD1,DRD5:::bin::D;ADA2A:::inh::D;5HT1D:::bin::D;5HT3A:::bin::D;5HT2C:::ant::D;HRH1:::ant::D;ADA2B;DRD2;ADA1B:::ant::D;ADA1A:::ant::D;5HT1A:::ant::D;5HT2A:::ago::D;SC6A3:::inh::D;SC6A2:::inh::D;SC6A4:::inh::D|CP2C9:::sub::D;CP2CJ:::sub::D;CP2D6:::sub::D|MDR1:::sub::D|
Nitroglycerin|ok_inv|ANPRA:::ago::D|ALDH2:::sub::D||
Rocuronium|ok|5HT3A:::ant::D;ACM2:::ant::D;ACHA2:::ant::D||SO1A2:::sub::D;S22A1:::sub::D|
Thiabendazole|ok_vet|MAP1::ECOLI::6.33:C;RAB9A::::5.6:C;HIF1A::::5.6:C;MAP11::::5.47:C;NPC1::::5.45:C;SMN::::5.2:C;CP2CJ::::5.1:C;P53::::5.:C;CP2D6::::5.:C;FRDA::ECOLI:inh::D|CP1A2:::inh:6.9:DC;CP1A1:::ind::D||
Nateglinide|ok_inv|S22A6::RAT::5.04:C;PPARG:::ago::D;ABCC8:::inh::D|CP2D6:::sub::D;UD19:::sub::D;PGH1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D|S22A6:::inh::D;S15A2:::inh::D;S15A1:::inh::D;MOT1:::sub::D;MRP4:::sub::D|A1AG1;ALBU
Atracurium_besylate|ok|ACHA2:::ant::D|||
Pralidoxime|ok_vet|TSHR::::6.2:C;CHLE:::act::D;ACES:::act::D|||
Risperidone|ok_inv|5HT2A:::ant:10.:DC;5HT2B::RAT::9.85:C;5HT2A::RAT::9.82:C;ADA1A::RAT::9.4:C;DRD2:::ant:9.36:DC;DRD2::RAT::9.27:C;ADA1A:::ant:9.16:DC;ADA1B::RAT::9.13:C;5HT7R::::9.:DC;ADA2C:::ago:8.86:DC;5HT7R::RAT::8.85:C;5HT2B::MOUSE::8.82:C;ADA2A:::ant:8.74:DC;HRH1:::ant:8.59:DC;ADA1D::::8.31:C;DRD4:::ant:8.21:DC;5HT2C:::ant:8.19:DC;DRD3:::ant:8.17:DC;ADA2C::RAT::8.1:C;HRH1::CAVPO::8.1:C;DRD3::RAT::8.01:C;5HT1B::::8.:C;ADA1B:::ant:8.:DC;ADA2B:::duo:7.92:DC;H10::::7.85:C;5HT2C::RAT::7.84:C;5HT2B::::7.82:C;DRD1:::ant:7.68:DC;5HT1A:::ant:7.68:DC;DRD1::RAT::7.66:C;DRD2::MOUSE::7.64:C;ADA2A::RAT::7.6:C;HRH1::RAT::7.1:C;5HT1A::RAT::6.89:C;KCNH2::::6.83:C;5HT6R::::6.65:C;GLRA1::::6.49:C;5HT1B::RAT::6.47:C;5HT1A::MOUSE::6.37:C;5HT1D:::ant:6.:DC;5HT5A::::6.:C;DRD5::::6.:C;SC6A4::::6.:C;HRH2::::5.84:C;CP2CJ::::5.8:C;S47A1::::5.8:C;ACM1::::5.55:C;SGMR1::::5.37:C;ACM3::::5.2:C;TSHR::::5.1:C|CP2D6:::inh:5.5:DC;CP3A4:::sub::D|MDR1:::sub::D|
Naftifine|ok|ERG2::YEAST::6.51:C;SGMR1::::6.06:C;EBP::::5.82:C;ERG1:::inh::D|||
Esomeprazole|ok_inv|ATP4A:::inh::D;DDAH1|CP2CJ:::inh::D;CP3A4:::sub::D|MDR1:::inh::D;S22A8:::inh::D|
Meclizine|ok|HEPS::::5.69:C;NR1I3:::ANT::D;HRH1:::ant::D|CP2D6:::sub::D||ALBU:::bin::D
Pentamidine|ok_inv|ACM4::::6.66:C;AOC1::::6.54:C;S47A1::::6.39:C;5HT2A::::6.33:C;ADA1A::RAT::6.31:C;ADA2A::::6.29:C;ACM2::::6.29:C;ADA1B::RAT::6.27:C;NMDZ1::::6.14:C;AOFA::::6.1:C;S100B::::6.:C;ST14::::5.94:C;S22A2::::5.92:C;NMDZ1::RAT::5.88:C;DRD3::::5.87:C;5HT2C::::5.77:C;SAT1::::5.7:C;ACM5::::5.68:C;SC6A2::::5.66:C;ACRO::PIG::5.64:C;SC6A3::::5.6:C;S47A2::::5.57:C;S22A3::::5.02:C;TRDMT;DNA:::itc::D|CP4AB:::sub::D;CP3A5:::sub::D;CP2D6:::sub::D;CP1A1:::sub::D;CP2CJ:::sub::D||
Hetacillin|ok_vet_out|PBP2A::STRR6:inh::D;PBP1B::STRR6:inh::D;PBP3::STREE:inh::D;PBPA::STRR6:inh::D;PBP2::STRR6:inh::D|||
Riluzole|ok_inv|SC6A2::::5.76:C;SCN2A::::5.66:C;RORG::MOUSE::5.55:C;PTR1::LEIMA::5.4:C;SCN2A::RAT::5.33:C;LYAG::::5.25:C;LMNA::::5.15:C;XCT:::ind::D;SCN5A:::inh::D|CP1A2:::sub:6.5:DC;CP1A1:::sub::D|ABCG2:::sub::D|
Hydrocortisone|ok_vet|GCR:::ago:7.92:DC;NFKB1::::7.85:C;GCR::MOUSE::7.37:C;HIF1A::::6.7:C;ACM1::RAT::6.6:C;TAU::::5.35:C;ANXA1:::ago::D|CP2CJ:::ind::D;CP2C9:::ind::D;CP2B6:::ind::D;CP1B1:::ind::D;CP2A6:::ind::D;DHI1:::sub::D;DHI2:::sub::D;S5A2:::sub::D;AK1D1:::sub::D;CP2C8:::ind::D;C11B2:::sub::D;C11B1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub_ind::D|S22A8:::sub::D;SO1A2:::inh::D;MDR1:::sub_ind::D|CBG:::bin:7.88:DC;SHBG:::bin:6.2:DC
Mannitol|ok_inv||O08355:::sub::D|MDR1:::sub::D|
Gadobenic_acid|ok_inv||||ALBU:::bin::D
Zileuton|ok_out|LOX5::RAT::6.85:C;LOX5::MOUSE::6.72:C;LMNA::::6.65:C;LOX5:::inh:6.52:DC;LT4R1::::6.38:C;AL5AP::::6.24:C;HYES::::6.23:C;LKHA4::::6.07:C|UD19:::sub::D;PGH1:::sub::D;CP3A4:::sub::D;CP1A2:::sub::D;CP2C9:::sub::D||ALBU
Modafinil|ok_inv|LMNA::::8.74:C;DRD2::::8.68:C;SC6A3:::inh:6.19:DC;SC6A3::RAT::5.6:C;ADA1B:::pag::D|CP3A5:::duo::D;CP2C9:::duo::D;CP2B6:::duo::D;CP1A2:::ind::D;CP3A4:::sub_ind::D;CP2CJ:::inh::D||
Deferoxamine|ok_inv|A4;Aluminum:::chel::D;Iron:::chel::D|XDH:::inh::D||
Scopolamine|ok_inv|ACM1:::ant::D;SUIS:::inh::D;ACM2:::ant::D;ACM3:::ant::D;ACM4:::ant::D;ACM5:::ant::D;ACHA4;ACHB2||MDR1:::inh::D|
Carbinoxamine|ok|HRH1:::ant::D|||
Etodolac|ok_inv_vet|BLM::::6.65:C;PGH2:::inh:6.25:DC;PGH1:::inh:5.58:DC;CP3A4::::5.5:C;RXRA|UD2B7:::sub::D;UD110:::sub::D;UD13:::sub::D;UD19:::sub::D;CP2C9:::sub::D|S22A6:::inh::D|ALBU
Prilocaine|ok|SCN5A:::inh::D|||
Epinastine|ok_inv|HRH1::CAVPO::8.85:C;S47A1::::5.96:C;S22A2::::5.37:C;5HT7R:::ant::D;5HT2A:::ant::D;ADA2A;ADA1A;HRH2:::ant::D;HRH1:::ant::D|CP3A4:::sub::D;CP2D6:::inh::D;CP2B6:::sub::D|MDR1:::sub::D|
Tranylcypromine|ok_inv|AOFB:::inh:5.98:DC;AOFA:::inh:5.92:DC;5HT2C::::5.57:C;CP2B6::::5.16:C|CP2A6:::inh:7.1:DC;CP2CJ:::inh:5.51:DC;CP2E1:::inh::D;CP1A2:::inh::D;CP2C9:::inh::D;CP2D6:::inh::D||
Isoflurane|ok_vet|ACHB2:::ant::D;ACHA4:::ant::D;GABAR:::aga::D;CALM1;ATPD;KCNA1:::ind::D;GRIA1:::ant::D;GLRA1:::ago::D;AT2C1:::inh::D;GBRA1:::ago::D|NU1M:::inh::D;CP2B6:::duo::D;CP2E1:::sub::D||ALBU
Ethotoin|ok|NR1I2:::act::D;SCN5A:::inh::D|||THBG:::sub::D
Tretinoin|ok_inv_nutra|RARG:::ago:10.4:DC;RARA::::10.:DC;RORB::::9.82:C;RARB::::9.4:DC;RABP1::MOUSE::9.4:C;RXRA::::9.4:DC;RXRB:::ago:9.3:DC;RXRG:::ago:8.85:DC;RABP2::MOUSE::8.7:C;RARB::MOUSE::8.7:C;RARG::MOUSE::8.4:C;RARA::MOUSE::8.3:C;RXRG::MOUSE::8.22:C;BLM::::7.65:C;RORG::::6.7:C;RORA::::6.7:C;5HT2B::::6.64:C;HIF1A::::6.6:C;RXRB::MOUSE::6.51:C;RABP1::CHICK::6.43:C;MK01::::6.24:C;RXRA::MOUSE::6.:C;AA3R::::5.53:C;RORG::MOUSE::5.3:C;HPGDS;CP26C;CP26B;CP26A;PDK4;RET4;OBP2A;LCN1;TIG1:::ago::D;AL1A2;NR0B1;RAI3;AL1A1|CP4AB:::sub::D;CP1A1:::sub::D;CP2CI:::sub::D;CP2A6:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP2B6:::sub::D;CP3A7:::sub::D|RABP2:::sub::D;RABP1:::sub::D|ALBU
Hexachlorophene|ok_out|MK14::::7.06:C;MK01::::6.71:C;STRP::STRP1::6.69:C;AA3R::::6.44:C;LMNA::::6.35:C;PGH2::::6.19:C;EGFR::::6.13:C;HS90A::::6.11:C;AA2AR::::6.04:C;ADA2C::::5.99:C;CP2CJ::::5.91:C;CP1A2::::5.88:C;NK2R::::5.86:C;DNAB::MYCTU::5.74:C;ADA2A::::5.69:C;ESR1::::5.67:DC;SC6A4::::5.64:C;5HT2C::::5.62:C;LCK::::5.61:C;MK03::::5.6:C;ACES::::5.52:C;THAS::::5.51:C;RORG::MOUSE::5.5:C;ANDR::RAT::5.48:C;ERBB2::::5.48:C;PAX8::::5.48:C;FYN::::5.46:C;5HT2B::::5.44:C;CAN2::PIG::5.43:C;LOX15::::5.3:C;TERA::::5.26:C;HD::::5.25:C;RECA::MYCTU::5.14:C;TAU::::5.1:C;HCD2::::5.1:C;NPY1R::::5.01:C;TSHR::::5.:C;DHE3:::inh::D;DHSD:::inh::D;DLD::ECOLI:inh::D|||
Dolasetron|ok_inv|KCNH2::::5.23:C;5HT3A:::ant::D|CP2C9:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D||
Clopidogrel|ok|SC6A4::::6.52:C;P2Y12:::ant::D|CP2B6:::inh:6.3:DC;EST1:::sub::D;CP2C8:::inh::D;CP1A2:::sub::D;CP2C9:::inh::D;CP2CJ:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|S22A2:::inh::D;S22A1:::inh::D;MDR1:::sub::D|
Tetracycline|ok_vet|PTN7::::5.08:C;PADI4;Multidrug_translocase_MdfA::ECOLX:::D;PRIO:::inh::D;16S_ribosomal_RNA::Gut_flora:inh::D;RS19::ECOLI:inh::D;RS8::ECOLI:inh::D;RS3::ECOLI:inh::D;RS14::ECOLI:inh::D;RS7::ECOLI:inh::D|CP3A4:::inh::D|SO2B1:::inh::D;S22A7:::inh::D;S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D|ALBU
Meropenem|ok_inv|STRP::STRP1::6.9:C;DACB::ECOLI:inh::D|BLO10::PSEAI:sub::D||
Potassium_chloride|ok_out|||S12A4:::sub::DC;S12A7:::sub::DC;S12A6:::sub::DC;S12A5:::sub::DC;S12A1:::sub::DC;S12A2:::sub::DC|
Irinotecan|ok_inv|ACES::TETCF::7.58:C;ACES::::7.3:C;ACM4::::6.66:C;ADA2C::::6.34:C;S47A1::::5.68:C;S22A2::::5.57:C;MMP1::::5.22:C;S47A2::::5.1:C;TOP1M:::inh::D;TOP1:::inh::D|CHLE:::sub::D;EST2:::sub::D;EST1:::sub::D;UD19:::sub::D;UD11:::sub::D;CP3A7:::sub::D;CP2B6:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|MRP2:::sub::D;MDR1:::sub::D;ABCG2:::sub::D;MRP1:::sub::D;SO1B1:::inh::D;S22A3:::inh::D|ALBU:::sub::D
Methimazole|ok|LMNA::::8.7:C;PERL::BOVIN::5.08:C;PERT:::inh::D|FMO3:::sub::D;CP3A4:::inh::D;CP2E1:::inh::D;CP2D6:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D;CP2B6:::inh::D;CP2A6:::inh::D;CP1A2:::inh::D||
Mometasone|ok_vet|GCR:::ago::D;PRGR:::ago::D|CP2C8:::inh::D;CP3A4:::sub_ind::D;CP3A5:::ind::D||
Metyrosine|ok|IMPA1::RAT::5.4:C;BLM::::5.25:C;TY3H:::bin::D|||
Clavulanic_acid|ok_vet|AMPC::ECOLI::7.82:C;BLA1::ECOLX::7.55:C;BLAT::ECOLX::7.53:C;BLAC::STAAU::7.1:C;BLA1::KLEPN::6.77:C;AMPC::PSEAE::6.1:C;BLO1::ECOLX::5.49:C|Bacterial_beta_lactamase_enzymes::UNK:inh::DC|SC5A1:::ind::D|
Olopatadine|ok|HRH1:::ant::D;HRH2:::ant::D;HRH3:::ant::D;S10A1:::ant::D;S10AC:::ant::D;S100B;S10AD;S10A2:::ant::D|CP3A4:::sub::D;FMO1:::sub::D;FMO3:::sub::D|MDR1:::sub::D|ALBU:::bin::D
Hydrocortamate|ok|GCR:::ago::D|CP3A4:::ind::D||
Alprostadil|ok_inv|PI2R::::8.74:C;PE2R4::MOUSE::8.6:C;PE2R2::MOUSE::8.59:C;PE2R3::MOUSE::8.3:C;PE2R1::MOUSE::8.22:C;SO2B1::RAT::7.45:C;PD2R2:::ago::D;PE2R1:::ago::D;PE2R2:::ago::D||S22A6:::inh::D;SO2A1:::sub::D;MRP4:::sub::D;SO3A1:::inh::D;SO2B1:::inh::D;MRP5:::inh::D|
Clidinium|ok|ACM1:::ant::D|||
Malathion|ok_inv|CP3A4::::6.:C;HCD2::::5.4:C;AL1A1::::5.25:C;CHLE:::inh::D|CP2B6:::sub::D;CP1A2:::sub::D||
Etoposide|ok|NCOA3::::6.43:C;LMP1::EBVB9::6.4:C;TOP2A:::inh:6.09:DC;NCOA1::::5.94:C;LOX15::RABIT::5.5:C;SO1B3::::5.38:C;TOP2B:::inh::D|PGH1:::sub::D;PGH2:::sub::D;GSTP1:::sub::D;GSTT1:::sub::D;UD11:::sub::D;CP3A5:::sub::D;CP2E1:::sub::D;CP1A2:::sub::D;CP3A4:::duo::D|ABCG2:::sub::D;MRP2:::inh::D;MRP7:::inh::D;MRP1:::inh::D;MDR1:::inh::D;MRP6:::inh::D;MRP3:::inh::D|
Hydroflumethiazide|ok_inv|LMNA::::6.:C;KCMA1;AT1A1;CAH12:::inh::D;CAH9:::inh::D;CAH4:::inh::D;CAH2:::inh::D;CAH1:::inh::D;S12A1:::inh::D|||
Tirofiban|ok|ITB3:::ant:9.43:DC;ITA2B:::ant::D|||
Oxcarbazepine|ok|SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A,SCN1B,SCN2B,SCN3B,SCN4B:::inh::D|CP3A5:::duo::D;CP3A4:::duo::D;CP2CJ:::inh::D;CBR3:::sub::D;CBR1:::sub::D;AK1C4:::sub::D;AK1C3:::sub::D;AK1C2:::sub::D;AK1C1:::sub::D|MDR1:::sub::D|ALBU:::sub::D
Propiomazine|ok|HRH1:::ant::D;5HT2A:::ant::D;5HT2C:::ant::D;DRD2:::ant::D;DRD1:::ant::D;DRD4:::ant::D;ADA1A:::ant::D;ADA1B:::ant::D;ADA1D:::ant::D;ACM3:::ant::D;ACM5:::ant::D;ACM2:::ant::D;ACM4:::ant::D;ACM1:::ant::D|||
Roxithromycin|ok_out|ADA1B::RAT::6.26:C;MDR1;RL10::SHIFL:inh::D|CP2B6:::inh::D;CP3A4:::inh::D||
Nalidixic_acid|ok_inv|LMNA::::6.9:C;RORG::MOUSE::5.55:C;DNA|CP1A2:::inh::D;T23O:::inh::D|S22A6:::inh::D|
Phenelzine|ok|NFKB1::::8.:C;AOC3:::inh:7.7:DC;AOFA::RAT::7.52:C;AOFB::RAT::7.12:C;TSHR::::6.9:C;CP2C9::::6.8:C;LMNA::::6.3:C;CP1A2::::6.:C;Glutamic_acid_decarboxylase:::inh::D;ALAT2:::inh::D;ALAT1:::inh::D;GABT:::inh::D|AOFB:::sub:7.03:DC;AOFA:::sub:6.84:DC;CP2CJ:::inh:6.5:DC;CP2D6:::inh:6.:DC;CP2C8:::inh:5.92:DC;CP3A4,CP343,CP3A5,CP3A7:::inh:5.7,,,:DC;CP3A4:::inh:5.7:DC;CP3A7:::inh::D;CP3A5:::inh::D;CP2E1:::ind::D||
Propantheline|ok|ACM1::RAT::9.:C;CP2D6::::5.9:C;TSHR::::5.1:C;ACM1:::ant::D|||
Estradiol|ok_inv_vet|ESR1:::ago:11.:DC;ESR2:::ago:11.:DC;ESR2::RAT::9.85:C;GPER1::::9.52:DC;ESR1::RAT::9.45:C;SMN::::8.85:C;ESR1::MOUSE::8.66:C;ESR2::MOUSE::8.64:C;ERR2::::8.49:C;ERR1::::8.44:C;ANDR::::7.72:C;BLM::::7.65:C;AOXA::::7.1:C;ANDR::RAT::6.63:C;S22A3::RAT::5.96:C;ST1A1::::5.92:C;TAU::::5.7:C;AOXA::RAT::5.52:C;LMNA::::5.45:C;CP2B6::::5.39:C;SO1A1::RAT::5.33:C;SC6A4::::5.24:C;CBG::::5.:C;ERR3:::lig::D;DHB2;BECN1;ATP6;NCOA2;ACHA4;NR1I2|CP3A4:::sub_ind:6.:DC;CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D;UD11:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP1A2:::inh::D|S22A3:::inh:5.54:DC;S22A1:::inh:5.24:DC;SO4A1;SO1C1;SO1B3;S22A8:::sub::D;MDR1:::sub::D;SO1B1:::inh::D;ABCG2:::duo::D;S22AB:::inh::D;MRP7:::inh::D;SO1A2:::inh::D;SO2B1:::inh::D;S22A2:::inh::D|SHBG::::8.83:DC;FABPI;ALBU
Mefenamic_acid|ok|TYDP1::::7.95:C;PGH1:::inh:6.94:DC;AK1C2::::6.66:C;AK1C3::::6.52:C;PGH2:::inh:6.22:DC;AK1C1::::6.09:C;AK1BA::::5.8:C;CP1A2::::5.3:C;ACES::TETCF::5.21:C;HIF1A::::5.:C;CP3A4::::5.:C|CP2C9:::sub:5.1:DC;UD19:::inh::D;CP2C8:::inh::D||ALBU
Cryptenamine|ok|ACM2:::ant::D;ACM1:::ant::D;ACM3:::ant::D;ACM4:::ant::D;ACM5:::ant::D|||
Acyclovir|ok|BLM::::6.3:C;RECQ1::::6.1:C;DPOL::VZVD:inh::D;DPOL::HHV11:inh::D;KITH::HHV11:pot::D|PURA1,PURA2:::sub::D;PCKGM,PCKGC:::sub::D;SUCB1,SUCA,SUCB2:::sub::D;PGK1,PGK2:::sub::D;KCRB,KCRM,KCRS,KCRU:::sub::D;KPYR,KPYM:::sub::D;NDKA,NDKB:::sub::D;KGUA:::sub::D;KITH::HHV1:sub::D|S47A2:::sub::D;S47A1:::sub::D;NTCP2:::sub::D;S22A8:::inh::D;S22A6:::inh::D;S22A1:::inh::D|ALBU:::bin::D
Naproxen|ok_vet|PGH2::RAT::7.22:C;PGH1::SHEEP::6.74:C;PGH1:::inh:6.68:DC;AK1C3::::6.32:C;TSHR::::6.1:C;LIPS::RAT::5.92:C;S22A6::RAT::5.7:C;PGH2:::inh:5.6:DC;PAB::FINMA:::D|CP1A2:::sub:5.:DC;UD110:::sub::D;UD19:::sub::D;UD18:::sub::D;UD17:::sub::D;UD16:::sub::D;UD13:::sub::D;UD2B7:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D|S22A6:::inh:5.24:DC;S22A8;MDR1:::inh::D;ABCBB:::sub::D;SO1A2:::inh::D|ALBU
Gadopentetic_acid|ok|6PGD:::inh::D|||
Perindopril|ok|ACE:::inh:8.82:DC;AMPC::ECOLI::5.35:C;SFRP4:::inh::D|CHLE:::inh::D|S15A2:::sub::D;S15A1:::sub::D|
Uracil_mustard|ok|DNA:::itc::D|||
Tripelennamine|ok_vet|HRH1:::ant:7.4:DC|CP2D6:::inh::D||
Haloprogin|ok_out|AA3R::::6.9:C;DRD3::::6.78:C;ADA2B::::6.6:C;DRD1::::6.55:C;SC6A4::::6.37:C;OPRK::::6.34:C;ADA2A::::6.34:C;NK2R::::6.31:C;GALE::::6.3:C;ADA2C::::6.23:C;5HT2A::::6.16:C;5HT2C::::5.87:C;SC6A3::::5.81:C;5HT6R::::5.73:C;SC6A2::::5.56:C;RORG::MOUSE::5.25:C;NR1I2::::5.:C|||
Primidone|ok_vet|TSHR::::5.2:C;GABAR:::aga::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|UD11:::ind::D;CP1A2:::ind::D;CP3A4:::ind::D;CP2C9:::sub_ind::D;CP2CJ:::sub_ind::D||
Sulfasalazine|ok|LMNA::::7.5:C;HIF1A::::6.65:C;TSHR::::5.8:C;CAH1::::5.52:C;CAH2::::5.35:C;MK01::::5.2:C;PA21B:::ant::D;THAS:::ant::D;THIL:::inh::D;XCT:::inh::D;IKKB:::inh::D;IKKA:::inh::D;PPARG:::ago::D;PGH1:::inh::D;PGH2:::inh::D;LOX5:::inh::D||SO1B1:::inh:6.28:DC;SO2B1:::inh:5.52:DC;SO1B3:::inh::D;PCFT:::inh::D;MRP2:::sub::D;ABCG2:::inh::D|
Candesartan_cilexetil|ok|AGTR1::RABIT::6.7:C;SO1B1::::6.4:C;SO1B3::::5.72:C;POLK::::5.25:C;POLI::::5.21:C;CYSP::TRYCR::5.2:C;AGTR1:::ant::D|PGH1:::sub::D;UD13:::sub::D;CP2C8:::inh::D;CP2C9:::sub::D|MDR1:::inh::D|
Tolazoline|ok_vet|LMNA::::6.75:C;ADA2C::RAT::6.74:C;TAAR1::::5.79:C;ADA1B::RAT::5.68:C;ADA1A:::ant:5.41:DC;CP1A2::::5.:C;ADA2B:::bin::D;ADA2C:::bin::D;HRH2:::ago::D;HRH1:::ago::D;ADA2A:::ant::D|||
Gentamicin|ok_vet|DYR;NADE::BACSU:::D;LRP2;16S_ribosomal_RNA::Gut_flora:cov::D;RS12::ECOLI:cov::D||S22A6:::inh::D|
Tazarotene|ok_inv|RARB:::ago:9.1:DC;RARG:::ago:7.4:DC;RARA:::ago:7.2:DC;RXRB:::ago::D|CP2C8:::sub::D||
Fenoldopam|ok|DRD1::RAT::8.91:C;DRD2::RAT::7.88:C;DRD1:::ago:7.55:DC;AA2BR::RAT::7.45:C;ADA1A:::inh:6.82:DC;DRD2::BOVIN::6.1:C;DRD2::::6.09:C;KDM4E::::5.72:C;DRD2:S197A:RAT::5.72:C;DRD2:S194A:RAT::5.57:C;ADA1D:::inh::D;ADA1B:::inh::D;ADA2A:::ant::D;ADA2C:::ant::D;ADA2B:::ant::D;DRD5:::ago::D|||
Halazepam|ok_ill_out|GABAR:::aga::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRA5:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|||
Alfentanil|ok_ill|OPRM::RAT::8.09:C;SGMR1::RAT::8.09:C;OPRM::CAVPO::7.82:C;OPRM:::ago::D|CP3A5:::sub::D;CP3A7:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|ALBU;A1AG1
Colistin|ok|MC3R::::6.77:C;MC5R::::6.6:C;MC4R::::6.09:C;FYN::::6.02:C;EGFR::::5.82:C;ERBB2::::5.65:C;Bacterial_outer_membrane::Bacteria:destbz::D|||
Dicyclomine|ok|ACM4::::9.39:C;ACM1:::ant:9.08:DC;ACM3::::9.03:C;ACM5::::8.77:C;SGMR1::::8.69:C;ACM1::RAT::8.61:C;ACM2:::ant:7.8:DC;ACM2::RAT::7.33:C;5HT2A::::7.16:C;LMNA::::7.15:C;5HT2C::::6.61:C;DRD3::::6.39:C;5HT2B::::6.08:C;5HT6R::::5.85:C;HRH2::::5.8:C;CP3A4::::5.6:C;CP1A2::::5.4:C;CP2D6::::5.3:C;TPO::::5.:C|||
Minaprine|ok|IMPA1::RAT::8.6:C;ACM1::RAT::5.22:C;CP3A4::::5.:C;CP1A2::::5.:C;ACM1:::ago::D;DRD2:::ago::D;DRD1:::ago::D;SC6A4:::inh::D;ACES:::inh::D;5HT2C:::ant::D;5HT2A:::ant::D;5HT2B:::ant::D;AOFA:::inh::D|CP2D6:::sub:5.1:DC||
Pentoxifylline|ok_inv|IMPA1::RAT::7.6:C;ACM1::RAT::7.15:C;AA2BR::::5.29:C;LMNA::::5.25:C;ACES::::5.18:C;5NTD:::inh::D;AA2AR:::ant::D;PDE4A:::inh::D;PDE5A:::inh::D;AA1R:::ant::D;PDE4B:::inh::D|CP1A2:::sub::D||
Proparacaine|ok_vet|SGMR1::::7.:C;CP3A4::::5.9:C;AOFA::::5.75:C;SCN1A::::5.72:C;LEF::BACAN::5.5:C;CP1A2::::5.3:C;CP2D6::::5.2:C;SCNAA:::inh::D|||
Indapamide|ok|CAH7::::9.64:C;CAH12::::8.:C;CAH13::MOUSE::7.89:C;CAH9::::7.44:C;CAH13::::7.:C;CAH2::::6.7:C;CAH4::::6.67:C;CAH6::::6.6:C;CAH5B::::6.56:C;CAH5A::::6.05:C;LOX15::RABIT::5.53:C;CAH14::::5.31:C;LYAG::::5.2:C;CAH1::::5.:C;S12A3:::inh::D|CP3A4:::sub::D||
Tropicamide|ok_inv|BLM::::8.46:C;ACM4:::ant:8.46:DC;ACM3:::ant:7.52:DC;ACM2:::ant:7.43:DC;ACM5::::7.19:C;ACM1:::ant:7.17:DC;END4::ECOLI::6.15:C;CP2CJ::::6.:C;CP2C9::::6.:C;TAU::::5.45:C|||
Biperiden|ok_inv|ACM1:::ant::D;ACHA2:::ant::D|CP2D6:::inh::D||
Ribavirin|ok|LMNA::::8.4:C;ACM1::RAT::7.3:C;CP3A4::::6.1:C;POLG::DEN2P:::D;ENPP1:::inh::D;5NTC:::ind::D;RDRP::I56A0:inh::D;L::PI2HT:ant::D;IMDH2;IMDH1:::inh::D|ADK:::act::D|S29A1:::sub::D;S28A3:::sub::D|
Phenylbutazone|ok_vet|LMNA::::8.:C;NPSR1::::6.5:C;AL1A1::::5.95:C;PGH1:::inh:5.52:DC;HCD2::::5.5:C;FPR1::::5.28:C;PTGIS:::inh::D;PGH2:::inh::D|CP3A4:::ind::D;CP2C9:::inh::D|S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D|
Fentanyl|ok_ill_inv_vet|SGMR1::RAT::8.94:C;OPRM:::ago:8.89:DC;OPRM::RAT::8.82:C;OPRM::CAVPO::8.51:C;OPRD::MOUSE::8.46:C;OPRM::MOUSE::8.23:C;OPRD:::ago:6.73:DC;OPRK:::ago:6.71:DC;OPRK::CAVPO::6.71:C;OPRD::RAT::6.4:C;KCNH2::::5.74:C;AOFA::::5.26:C|CP3A7:::sub::D;CP3A4:::sub::D|MDR1:::inh:5.19:DC|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Meloxicam|ok_vet|PGH2::MOUSE::6.82:C;PGH2:::inh:6.8:DC;PGH1::SHEEP::6.:C;PGH1:::inh:5.88:DC;PGH2::SHEEP::5.86:C|CP2C8:::inh::D;6PGD:::inh::D;CP3A4:::sub::D;CP2C9:::sub::D|MRP4:::sub::D|
Sodium_lauryl_sulfate|ok|LEF::BACAN::7.:C|||ALBU:::bin::D
Orciprenaline|ok|ADRB2:::ago:6.3:DC;RORG::MOUSE::5.25:C;ADRB2::BOVIN::5.04:C|||
Rosoxacin|ok_inv|PARC::ECOLI:inh::D;GYRB::ECOLI:inh::D|CP1A2:::inh::D||
Propofol|ok_inv_vet|LMNA::::5.95:C;GBRA1::::5.7:C;5HT2B::::5.46:C;PGH1::::5.42:C;GBRP::RAT::5.4:C;5HT2C::::5.22:C;LOX15::RABIT::5.12:C;SC6A2::::5.03:C;GABAR:::aga::D;SCN2A:::inh::D;SCN4A:::inh::D;GBRB3:::pot::D;GBRB2:::pot::D|CP1A2:::inh:5.:DC;UD16:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP2CI:::sub::D;CP1A1:::inh::D;CP1B1:::inh::D;CP2E1:::inh::D;FAAH1:::sub::D;UD11:::inh::D;UD19:::sub::D;UD18:::sub::D;CP2B6:::sub::D;CP2C9:::sub::D||ALBU
Acetazolamide|ok_vet|CAH9::::10.22:C;CAH2:::inh:9.1:DC;CAH5B::::8.74:C;CAH7:::inh:8.6:DC;CAH12:::inh:8.6:DC;CAH3:::inh:8.51:DC;CAH14:::inh:8.24:DC;CAH13::::8.24:C;MTCA2::MYCTU::8.05:C;CAH6::::7.96:C;CAH4:::inh:7.96:DC;CAH1:::inh:7.92:DC;CAH2::BOVIN::7.8:C;CAH7::MOUSE::7.8:C;CAH13::MOUSE::7.77:C;CYNT::HELPY::7.7:C;CAHX::FLABI::7.57:C;CAN::CANAL::7.4:C;CAH5A::::7.22:C;CAH::METTE::7.22:C;CAH4::BOVIN::7.15:C;CAH15::MOUSE::7.14:C;CAN::YEAST::7.09:C;MTCA1::MYCTU::6.6:C;THB::::5.75:C;MEN1::::5.05:C;AQP1:::inh::D|CP3A4:::inh::D|S22A6:::inh::D|
Tadalafil|ok_inv|PDE5A:::inh:8.92:DC;PDE5A::BOVIN::8.48:C;PDE5A::RAT::8.3:C;PDE11:::inh:8.:DC;CNCG::::6.01:C;PDE6A::BOVIN::5.52:C;MK01::::5.4:C;PDE6B::BOVIN::5.29:C;PDE4A::::5.04:C|CP3A5:::sub::D;CP3A4:::sub::D||
Carprofen|ok_vet_out|PGH2:::inh:7.:DC;PGH1:::inh::D||S22A6:::inh::D|
Disulfiram|ok|TAU::::7.6:C;LOX15::::7.2:C;MTOR::::7.18:C;LMNA::::7.05:C;AL1A1::::7.05:C;HCD2::::6.8:C;AA3R::::6.7:C;RORG::MOUSE::6.6:C;DRD3::::6.43:C;TPO::::6.4:C;CP2C9::::6.4:C;HD::::6.1:C;CP2CJ::::6.1:C;CCR2::::6.02:C;DRD1::::5.97:C;DRD4::::5.96:C;MGLL::::5.9:C;OPRM::::5.85:C;ADA2B::::5.83:C;MK03::::5.82:C;CP1A2::::5.8:C;PLIN5::::5.79:C;ADA2A::::5.74:C;LOX12::::5.7:C;FFP::BACIU::5.7:C;5HT1B::RAT::5.67:C;OPRK::::5.61:C;PGDH::::5.6:C;TRPA1::::5.52:C;SC6A3::::5.43:C;PTBP1::::5.4:C;LEF::BACAN::5.4:C;CXCR2::::5.38:C;CCR4::::5.36:C;CYSP::TRYCR::5.35:C;HS90A::::5.29:C;AGTR1::::5.18:C;ABHD5::::5.16:C;NFKB1::::5.15:C;5HT6R::::5.13:C;DRD2::::5.12:C;NPSR1::::5.1:C;DOPO:::inh::D;ALDH2:::inh::D|CP3A4:::sub:5.1:DC;CP3A5:::sub::D;CP2E1:::inh::D|ABCBB:::sub::D|
Ethynodiol_diacetate|ok|ANDR::RAT::5.68:C;AOFA::::5.37:C;ESR1:::ago::D;PRGR:::ago::D|CP3A4:::sub::D||
Enprofylline|ok_exp|BLM::::6.7:C;PGDH::::5.45:C;AA2BR:::ant:5.33:DC;HCD2::::5.2:C;AA2AR:::inh:5.14:DC;AA3R:::inh::D;AA1R:::inh::D;PDE4B:::inh::D;PDE4A:::inh::D|||
Levomenthol|ok|CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1A:::ant::D;OPRK:::ago::D;TRPV3:::ind::D;TRPA1:::ind::D;TRPM8:::ind::D|CP3A4:::sub::D||
Natamycin|ok|Ergosterol::CANAL:bin::D|CP3A4:::inh::D||
Cinoxacin|ok_out|LMNA::::8.3:C;BLM::::6.55:C;TSHR::::5.1:C;DNA:::itc::D;GYRA::HAEIN:inh::D|CP1A2:::inh::D|S22A6:::inh::D|
Fosfomycin|ok|MURA::ECOLI:inh:7.:DC|||
Diazepam|ok_ill_inv_vet|GBRG2::RAT::8.68:C;GBRP::RAT::8.54:C;GBRG1::RAT::8.3:C;GBRG2:::pot:8.18:DC;GBRA1:::pot:8.09:DC;GBRA2::BOVIN::8.:C;GBRB2:::pot:8.:DC;GBRA5::MOUSE::7.92:C;AA3R::::7.92:C;GBRA2::RAT::7.82:C;GBRA5:::pot:7.64:DC;CHLE::HORSE::7.37:C;TSPO::RAT::6.71:C;FABPL::RAT::6.27:C;AK1C2::::5.62:C;AK1C1::::5.25:C;GABAR:::aga::D;TSPO:::pot::D;GBRT:::pot::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRG3:::pot::D;GBRG1:::pot::D;GBRB3:::pot::D;GBRB1:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D|CP2E1:::inh::D;PGH1:::sub::D;CP2C8:::sub::D;CP2CI:::sub::D;CP2B6:::sub::D;CP2C9:::sub::D;CP2CJ:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::inh::D|MDR1:::sub::D|ALBU
Phenmetrazine|ok_ill|SC6A2:::inh::D;SC6A3:::inh::D|||
Trifluoperazine|ok_inv|DRD2::RAT::9.27:C;5HT2B::RAT::8.98:C;EBPL::::8.41:C;EBP::::8.1:C;SGMR1::::7.82:C;ADA1B::RAT::7.53:C;HCD2::::6.7:C;CP2D6::::6.5:C;5HT1A::RAT::6.39:C;ERG2::YEAST::6.3:C;CALM1:::inh:6.:DC;TAU::::5.9:C;PDR5::YEAST::5.85:C;CP2CJ::::5.7:C;CALM::BOVIN::5.47:C;SCN1A::::5.3:C;KCNH2::::5.29:C;BGLR::RAT::5.11:C;UBP1::::5.1:C;LYSC1::RAT::5.05:C;ACM1::RAT::5.:C;CP3A4::::5.:C;LEF::BACAN::5.:C;S10A4:::inh::D;TNNC1;ADA1A:::ant::D;CALY:::ant::D;DRD2:::ant::D|CP1A2:::sub:6.2:DC;UD14:::sub::D;XDH:::inh::D|MDR1:::inh:5.2:DC|
Phensuximide|ok|AMPC::ECOLI::5.25:C|||
Cefaclor|ok|STRP::STRP1::6.33:C;CTDS1::::5.14:C;PBPA::CLOPE:inh::D;PBP3::STREE:inh::D|PERM:::ind::D|ABCBB:::sub::D;S22A8:::inh::D;S15A2:::inh::D;S15A1:::inh::D|
Mifepristone|ok_inv|PRGR:::ant:10.68:DC;GCR:::ant:10.:DC;ANDR::::9.19:C;VP16::HHV11::9.15:C;GCR::RAT::8.85:C;GCR::MOUSE::8.66:C;PRGR::RAT::8.46:C;ANDR::RAT::8.25:C;LOX15::RABIT::6.26:C;MCR::::6.23:C;ESR2::::6.09:C;OPRM::::6.:C;FRIL::HORSE::5.7:C;ESR1::::5.3:C;LMNA::::5.25:C;OPRK::::5.09:C;RORG::MOUSE::5.05:C;NR1I2;KLK3|CP3A4:::duo:5.33:DC;CP2C9:::inh::D;CP2C8:::inh::D;CP2D6:::inh::D;CP3A5:::sub::D|SO1B3:::inh::D;SO1B1:::inh::D;ABCBB:::sub::D;MRP1:::inh::D;MDR1:::duo::D|
Brompheniramine|ok|SC6A4::RAT::6.52:C;KCNH2::::6.05:C;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;HRH1:::ant::D|||
Loperamide|ok|OPRM::RAT::9.8:C;OPRM:::ago:9.28:DC;OPRD::RAT::7.3:C;OPRM::CAVPO::7.24:C;OPRD:::ago:6.81:DC;SGMR1::::6.58:C;SCN1A::::6.57:C;DRD3::::6.34:C;ADA1B::RAT::6.27:C;SC6A4::::5.93:C;TSHR::::5.9:C;OPRK:::ago:5.9:DC;ADRB2::::5.68:C;ADA1A::RAT::5.6:C;5HT2B::::5.58:C;HRH2::::5.52:C;CALM::BOVIN::5.46:C;LMNA::::5.45:C;RORG::MOUSE::5.4:C;TIE2::::5.23:C;NR1I3;CALM1:::inh::D;COLI:::mod::D;CAC1A:::inh::D|CP2D6:::sub:7.8:DC;CP3A4:::inh:5.3:DC;CP2B6:::sub::D;CP2C8:::sub::D|MDR1:::sub:5.6:DC|
Progabide|exp|GBRA1:::ago::D;GABR1:::ago::D|||
Clocortolone|ok|GCR:::ago::D|||
Tolazamide|ok_inv|ACM1::RAT::7.95:C;END4::ECOLI::6.95:C;LOX15::RABIT::5.29:C;AGAL::::5.25:C;LOX12::::5.15:C;ABCC8,KCJ11:::inh::D|CP2C9:::sub::D||
Hydroxypropyl_cellulose|ok||||
Dobutamine|ok|ADA1A::RAT::7.35:C;ADA1D::::7.25:C;SC6A3::::6.91:C;ADA1B::RAT::6.73:C;SC6A2::::6.42:C;CAH15::MOUSE::6.41:C;CAH2::::6.32:C;LOX15::RABIT::6.22:C;CAH5A::::6.14:C;CAH5B::::6.05:C;SC6A4::::6.:C;ADRB2:::ago:5.98:DC;SGMR1::::5.98:C;ADRB1:::ago:5.95:DC;ADA2B::::5.87:C;DRD3::::5.77:C;CAH1::::5.72:C;FYN::::5.4:C;CAH7::::5.37:C;CAH12::::5.36:C;EGFR::::5.26:C;LCK::::5.26:C;CAH3::::5.13:C;CAH4::::5.05:C;CAH6::::5.02:C;CAH13::::5.02:C;CAH9::::5.01:C;ESR1;ADA1A,ADA1B,ADA1D:::ago:,,7.25:DC|COMT:::sub::D||
Oxazepam|ok|LMNA::::6.35:C;GABAR:::aga::D;GBRT:::pot::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|UD19:::sub::D;UD2B7:::sub::D;UDB15:::sub::D||
Donepezil|ok|ACES::RAT::8.77:C;ACES:::inh:8.7:DC;ACES::BOVIN::8.54:C;ACES::ELEEL::8.37:C;CLAT::RAT::8.28:C;ACES::MOUSE::8.05:C;ACES::TETCF::7.92:C;SGMR1::::7.84:C;CHLE:::ind:7.7:DC;HRH3::::6.46:C;CHLE::HORSE::6.27:C;KCNH2::::5.7:C;BACE1::::5.49:C;NMDA:::rdw::D;NFKB2,NFKB1:::inh::D;IL1B:::duo::D;TSG6:::inh::D;NOS1:::duo::D;5HT2A:::ind::D|CP2C9:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D|MDR1:::sub::D;ABCG2:::sub::D|
Nalbuphine|ok|OPRM:::ant:9.05:DC;OPRK:::ago:8.66:DC;OPRD:::ant:6.62:DC|||
Clofazimine|ok_inv|STRP::STRP1::5.91:C;CP2D6::::5.6:C;HIF1A::::5.6:C;MEN1::::5.5:C;MK01::::5.5:C;CYSP::TRYCR::5.22:C;CZCO::GEOKA:inh::D;DNA:::itc::D|CP3A4:::duo::D|MDR1:::inh:6.22:DC;ABCBB:::inh::DC|
Flurandrenolide|ok|GCR:::ago:8.69:DC;HIF1A::::8.2:C;NPSR1::::6.5:C|CP3A4:::sub::D||CBG:::bin::D
Cysteamine|ok_inv|CP3A4::::6.:C;NPY2R;SMS:::bin::D;Cystine:::cli::D|PERM:::sub::D||
Levamisole|ok_inv_vet_out|PPBT::BOVIN::5.74:C;ACH2::CAEEL:act::D;ACH7::CAEEL:act::D;ACH6::CAEEL:act::D;ACH5::CAEEL:act::D;PPBN:::inh::D;ACHA3:::ago::D|||
Methylphenobarbital|ok|LMNA::::6.35:C;NR1I2:::act::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2B6:::sub::D;CP2CJ:::sub::D||
Perphenazine|ok|DRD2:::ant:9.52:DC;5HT7R::::7.64:C;AOXA::::7.48:C;AOXA::RAT::6.13:C;PDR5::YEAST::5.85:C;KCNH2::::5.46:C;AOXA::MACFA::5.44:C;AOXA::MOUSE::5.21:C;END4::ECOLI::5.2:C;MTOR::::5.13:C;TAU::::5.05:C;P53::::5.:C;NPSR1::::5.:C;CALM1:::inh::D;DRD1:::ant::D|CP2D6:::inh:7.5:DC;CP1A2:::sub:6.5:DC;CP3A4:::sub:5.6:DC;CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP2CI:::sub::D||
Dacarbazine|ok_inv|MMP9::::6.25:C;6PGD:::inh::D;DPOA2;DNA:::cov::D|CP2E1:::sub::D;CP1A2:::sub::D;CP1A1:::sub::D||
Pseudoephedrine|ok|LEF::BACAN::7.9:C;TSHR::::6.9:C;LOX15::::6.4:C;HCD2::::6.2:C;CP2C9::::6.1:C;CP2CJ::::5.8:C;TPO::::5.5:C;LOX12::::5.5:C;KPYM::::5.1:C;GNAI1::::5.1:C;KPYK::LEIME::5.:C;IL2:::inh::D;ATF1,ATF2,ATF3,ATF4,ATF5,ATF6A,ATF7,JDP2,FOS,JUN:::inh::D;NFKB1:::inh::D;TNFA:::inh::D;NFAC1:::inh::D;ADRB1:::ago::D;ADRB2:::pag::D;SC6A4:::inh::D;ADA2A:::ago::D;ADA1A:::ago::D;SC6A3:::inh::D;SC6A2:::inh::D|AOFA:::inh::D||
Temozolomide|ok_inv|MEN1::::5.:C;DNA:::cov::D|||
Levorphanol|ok|OPRM:::ago:9.89:DC;OPRM::CAVPO::9.68:C;OPRM::MOUSE::9.52:C;SGMR1::MOUSE::8.72:C;OPRK:::ago:8.64:DC;OPRK::CAVPO::8.64:C;OPRD:::ago:8.54:DC;OPRK::MOUSE::8.:C;NMDZ1::RAT::5.92:C;NMDZ1::::5.6:C|||
Aminolevulinic_acid|ok|HEM2:::ind::D||S15A2:::inh::D;S15A1:::inh::D|
Chlorphenesin|ok_exp||CP19A:::ind::D;CP3A4:::ind::D;XDH:::inh::D;PGH2:::inh::D;CHLE:::ind::D||
Terbinafine|ok_inv_vet|LMNA::::7.8:C;ERG1:::inh:7.52:DC;SGMR1::::6.63:C;ADA2A::::5.67:C;SC6A2::::5.39:C;ERG1::CANAL:inh::D|CP2D6:::inh:6.7:DC;PGH1:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP3A4:::sub_ind::D;CP1A2:::sub::D;CP2C9:::sub::D|MDR2::TRIIM:sub::D|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Penicillamine|ok|TAU::::5.1:C;Copper:::chel::D||SO1B1:::sub::D|
Prednisolone|ok_vet|MCR::::9.54:C;GCR:::ago:9.28:DC;GCR::MOUSE::8.47:C;IL6::::8.38:C;ADA17::::7.83:C;GCR::RAT::7.71:C;GLNA::::7.49:C;GPBAR::::6.6:C;PRGR::::5.68:C;ANDR::::5.6:C;FABPL::RAT::5.58:C|CP3A4:::sub_ind::D|MDR1:::sub::D;SO1A2:::inh::D|CBG:::bin:7.51:DC;ALBU:::bin::D
Diflunisal|ok_inv|RORG::MOUSE::7.2:C;LMNA::::5.65:C;CAH2::::5.57:C;CAH1::::5.47:C;HIF1A::::5.3:C;AL1A1::::5.05:C;PGH1:::inh::D;PGH2:::inh::D|UD19:::inh::D;UD18:::sub::D|S22A6:::inh:6.07:DC|TTHY::::6.24:DC;ALBU::::5.91:DC;TTHY:V30M:::5.25:DC
Vardenafil|ok|PDE5A:::inh:9.7:DC;CNCG:::alo:9.:DC;PDE11::::6.89:C;PDE1A::::6.64:C;PDE9A::::6.34:C;PDE3A::::6.24:C;PDE10::::6.1:C;PDE7A::::5.72:C;PDE2A::::5.51:C;PDE4A::::5.42:C;CNRG:::alo::D|CP3A5:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|
Ranitidine|ok|HRH2:::ant::D;ACES:::inh::D|CP1A2:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D;ACES:::inh::D|S22A1:::inh::D;MDR1:::inh::D;S22A8:::sub::D;S22A2:::sub::D|
Tacrolimus|ok_inv|FKB1A:::inh:9.7:DC;FKB1B::::9.4:C;MTOR::::9.02:C;SF3B3::::7.96:C;PP2BA::::7.83:C;FKBP5::::7.1:C;NR1I2::::5.3:C|CP3A4:::sub:6.92:DC;CP3A5:::sub:6.85:DC|SO1B1:::inh:5.43:DC;ABCA5:::sub::D;MDR1:::duo::D|A1AG1:::sub::D;ALBU:::sub::D
Benzphetamine|ok_ill|VMAT2:::ind::D;ADA2A:::ago::D;ADA1A:::ago::D;SC6A3:::inh::D|CP3A4:::sub::D;CP2B6:::sub::D;NCPR:::sub::D||
Alprenolol|exp_out|ADRB2:::ant:9.53:DC;ADRB1:::ant:8.64:DC;ADRB2::BOVIN::8.53:C;ADRB3:::ant:7.12:DC;5HT1A::RAT::6.93:C;FDFT::RAT::5.38:C;5HT1A:::ant::D|CP2D6:::sub::D||
Ritodrine|ok_inv|ADRB2::RAT::7.62:C;ADRB3::RAT::6.72:C;ADRB2:::ago::D|6PGD:::inh::D||
Benzonatate|ok|CP3A4::::5.2:C;CYSP::TRYCR::5.1:C;AMPC::ECOLI::5.05:C;SCN5A:::ant::D|||
Dorzolamide|ok|CAH2:::inh:10.37:DC;CAH12::::8.52:C;CAH7::::8.46:C;CAN::CANAL::8.05:C;CAH6::::8.:C;CAH13::MOUSE::7.74:C;CAH13::::7.74:C;CAH14::::7.57:C;CAH5B::::7.48:C;CAH5A::::7.38:C;CAH4:::inh:7.37:DC;CAH4::BOVIN::7.37:C;CAH9::::7.28:C;CAH15::MOUSE::7.21:C;MTCA2::MYCTU::7.:C;CAN::YEAST::6.96:C;CAH::METTE::6.39:C;CAH1:::inh:6.3:DC;MTCA1::MYCTU::6.13:C;CYNT::HELPY::5.37:C;CAH3:::inh:5.1:DC|CP2C9:::sub::D||
Suprofen|ok_out|PGH1:::inh:6.25:DC;PGH2:::inh:5.56:DC;IMPA1::RAT::5.3:C;AMPC::ECOLI::5.2:C|CP2C9:::inh:5.43:DC;UD2B7:::sub::D;UD11:::sub::D||
Terbutaline|ok|ADRB2:::ago:5.6:DC;ADRB2::BOVIN::5.4:C;ADRB1:::ant::D;ADRB3:::ago::D|CHLE:::inh::D||
Conivaptan|ok_inv|V2R:::ant:9.44:DC;V1AR:::ant:9.37:DC|CP3A4:::inh::D||
Loteprednol_etabonate|ok|GCR:::ago::D|CP3A4:::sub::D;PON1:::sub::D||
Guaifenesin|ok_inv_vet|NMDA:::ant::D|||
Flupentixol|ok_out|DRD1::RAT::9.52:C;SGMR1::::8.65:C;DRD5::RAT::8.52:C;KCNK2::::5.7:C;UBP1::::5.15:C;FFP::BACIU::5.1:C;MEN1::::5.:C;ACM1:::ant::D;ADA1A:::ant::D;DRD1:::ant::D;5HT2A:::ant::D;DRD2:::ant::D|DDC:::ind::D|MDR1:::inh::D|
Eprosartan|ok|AGTRB::RAT::9.:C;AGTR2::RAT::9.:C;AGTR1:::ant:8.7:DC||MRP2:::ind::D|
Sirolimus|ok_inv|MTOR:::inh:10.:DC;FKB1B::::9.7:C;FKB1A::::9.7:DC;IF4E::::9.3:C;FKBP5::::8.52:C;PDCD4::::7.3:C;RORG::MOUSE::6.95:C;NR1I2::::6.05:C;CP2C9::::5.7:C;CP2CJ::::5.4:C;FGF2|CP3A4:::sub:5.7:DC;CP3A7:::sub::D;CP3A5:::sub::D|SO1B1:::inh:5.96:DC;MDR1:::duo:5.9:DC;S47A1|
Chlorhexidine|ok_vet_out|P53::::8.1:C;LMNA::::7.45:C;S22A1::::6.68:C;S22A2::::6.4:C;S22A3::::6.39:C;S47A2::::6.3:C;S47A1::::6.15:C;RAD52::::5.77:C;MC4R::::5.7:C;TYTR::TRYCR::5.7:C;UBE2N::::5.66:C;RORG::MOUSE::5.45:C;PAX8::::5.24:C;RCE1::YEAST::5.24:C;MMP2::::5.12:C;MMP9::::5.12:C;CP2CJ::::5.1:C;CP2D6::::5.1:C;HKDC1::::5.05:C;CAT4::PSEAE:inh::D;HNMT:::inh::D;Bacterial_outer_membrane::Bacteria:destbz::D|||
Emtricitabine|ok_inv|Reverse_transcriptase_RNaseH::9HIV1:inh::D|DCK:::sub::D|S47A1:::sub::D|ALBU:::bin::D
Chlorothiazide|ok_vet|LMNA::::6.05:C;NFKB1::::5.4:C;TSHR::::5.1:C;CP3A4::::5.:C;CAH2:::inh::D;CAH1:::inh::D;S12A3:::inh::D||S22A6:::inh::D|
Quinapril|ok_inv|ACE:::inh:8.08:DC;ACE::RABIT::6.96:C|EST1:::sub::D|S22A8:::sub::D;S15A2:::sub::D;S15A1:::sub::D|ALBU:::bin::D
Clomifene|ok_inv|ESR1:::duo::D;SHBG|CP17A:::inh::D|MDR1:::sub::D|
Isosorbide_dinitrate|ok_inv|AMPC::ECOLI::5.25:C;ANPRA:::ago::D|CP2E1:::inh::D||
Risedronic_acid|ok_inv|FPPS:::inh:9.44:DC;Hydroxylapatite:::ant::D|PGH2:::ind::D||
Pemirolast|ok_inv||||
Bumetanide|ok|HIF1A::::6.1:C;NPSR1::::5.5:C;S22A6::RAT::5.26:C;LMNA::::5.25:C;TSHR::::5.2:C;UBP2::::5.2:C;CFTR:::ant::D;S12A5:::inh::D;S12A4:::inh::D;S12A2:::inh::D;S12A1:::inh::D|PGH2:::ind::D|SO1A2:::sub::D;S22A7:::inh::D;S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D;NTCP:::inh::D|
Mechlorethamine|ok_inv|DNA:::itc::D|CHLE:::inh::D||
Granisetron|ok_inv|5HT3A:::ant::D|CP3A4:::sub::D;CP1A1:::sub::D||
Dienestrol|ok_inv|AMPC::ECOLI::6.5:C;LMNA::::5.7:C;CP3A4::::5.1:C;TAU::::5.05:C;HIF1A::::5.:C;SHBG;ESR1:::ago::D|||
Sulfapyridine|ok|FFP::BACIU::6.2:C;CYSP::TRYCR::5.6:C;DHP1::MYCFO:inh::D|CP2C9:::inh::D||
Oxybuprocaine|ok_inv|LEF::BACAN::6.8:C;CP1A2::::6.4:C;SCN1A::::5.54:C;CP2D6::::5.2:C;HIF1A::::5.:C;SCNAA:::inh::D|CHLE:::sub::D||
Iron_Dextran|ok_vet|HBB:::act::D;HBA:::act::D;FRIH;FRIL|||TRFE:::sub::D
Testolactone|ok_inv|CP19A:::inh::D|||
Benzylpenicilloyl_polylysine|ok|FCERG:::ago::D;FCERA:::ago::D|||
Rimexolone|ok|NR1I2::::6.4:C;NR1I2::RAT::6.17:C;AMPC::ECOLI::5.55:C;GCR:::ago::D|CP3A5:::ind::D;CP3A4:::sub_ind::D||CBG:::bin::D
Triazolam|ok_inv|GBRG2:::pot:9.23:DC;GBRA1:::pot:9.1:DC;GBRP::RAT::9.1:C;GBRA5:::pot:8.4:DC;RORG::MOUSE::6.1:C;GABAR:::aga::D;TSPO;GBRT:::pot::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRG3:::pot::D;GBRG1:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRA6:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D|CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D||
Ethanol|ok|TSHR::::7.5:C;L1CAM;KCNJ9;CCG2;5HT3C;5HT3D;5HT3B;5HT3E;S29A2;GBRD;GBRT;GBRP;GBRE;GBRG3;GBRG1;ACHB3;ACHA6;ACHA5;ACHA3;ACHB4;CAC1D;CAC1S;GBRB2;GBRB3;GBRB1;ACHA9;ACHA7;KCNJ5;S29A1;VCAM1;KCNJ6;KCNJ3;ACHB2;ACHA4;GRIA3;GRIA4;GRIA2;GBRA6;ACHA2;CCG1;GRIA1;GBRA3;GBRA4;GBRA5;CAC1C;ACH10;GBRA2;5HT3A;CACB1;GLRA2:::ago::D;GLRA1:::ago::D;NMD3A:::ant::D;GBRA1:::ago::D|AK1A1:::sub::D;ADH6:::sub::D;ADH7:::sub::D;ADH4:::sub::D;ADHX:::sub::D;ADH1G:::sub::D;ADH1B:::sub::D;ADH1A:::sub::D;CP4AB:::ind::D;CP3A4:::duo::D;CP2E1:::sub_ind::D;CP2CJ:::inh::D;CP2C9:::inh::D;CP2B6:::inh::D;CP1A2:::sub::D;CP1A1:::inh::D||
Remifentanil|ok|OPRK:::ago::D;OPRD:::ago::D;OPRM:::ago::D|||
Didanosine|ok|PNPH;Reverse_transcriptase_RNaseH::9HIV1:inh::D||S29A2;S29A1;S22A6:::sub::D|ALBU
Bitolterol|out|ADRB2|||
Methdilazine|ok|HRH1:::ant::D|||
Etacrynic_acid|ok_inv|CP2C9::::6.2:C;ALDR::RAT::5.94:C;LMNA::::5.5:C;GSTP1:::inh:5.47:DC;ABHD5::::5.38:C;PLIN5::::5.32:C;GSTA1::::5.3:C;HD::::5.25:C;LEF::BACAN::5.2:C;TAU::::5.05:C;LEF1;S12A1:::inh::D;AT1A1:::inh::D|GSTA2:::inh::D|S22A6:::inh::D|ALBU
Ondansetron|ok|5HT3A:::ant:10.1:DC;5HT3A::RAT::9.8:C;5HT3B::MOUSE::7.92:C;S47A1::::7.52:C;5HT3A::CAVPO::6.9:C;S47A2::::6.8:C;KCNH2::::6.4:C;5HT2B::::6.34:C;SGMR1::RAT::6.17:C;GASR::RAT::6.17:C;S22A2::::6.05:C;5HT4R::RAT::5.92:C;OPRM::RAT::5.54:C;5HT1B::RAT::5.43:C;5HT2C::RAT::5.3:C;5HT2B::RAT::5.:C;GBRP::RAT::5.:C;ACM1::RAT::5.:C;5HT1B;5HT1A;OPRM;5HT4R:::ago::D|CP2E1:::sub::D;CP2C9:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP2D6:::sub::D;CP1A2:::inh::D;CP3A4:::sub::D||
Bimatoprost|ok_inv|AK1C3::::5.3:C;PE2R3:::ago::D;PE2R1:::ago::D;PF2R:::ago::D|CP3A5:::sub::D;CP3A4:::sub::D||
Tiagabine|ok_inv|SC6A1:::inh:7.77:DC;SC6A1::MOUSE::7.43:C;SC6A1::RAT::7.15:C;S6A12::MOUSE::6.74:C|UD11:::sub::D;CP3A4:::sub::D||
Cocaine|ok_ill|SC6A4::RAT::9.3:C;KCNH2::::8.36:C;SC6A3::RAT::7.49:C;SC6A3:::inh:7.49:DC;SC6A4:::inh:7.35:DC;SC6A3::BOVIN::7.19:C;SC6A3::MACFA::7.02:C;SC6A2:::inh:6.97:DC;SGMR1::::5.05:DC;EST1;ACM2:::ant::D;ACM1:::ant::D;SCNAA:::inh::D;SCNBA:::inh::D;SCN5A:::inh::D|CHLE:::sub::D;CP2C8:::inh::D;CP2D6:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|S22A2:::inh::D|
Quinidine|ok_inv|TYDP1::::7.5:C;KCNH2:::inh:6.52:DC;CHLE::::5.91:C;KCND2::RAT::5.66:C;CP2DQ::RAT::5.55:C;SCN1A::::5.49:C;CAC1C::RAT::5.25:C;S22A1::RAT::5.22:C;CAC1C::::5.19:C;SCN5A:::inh:5.16:DC;KCNA5::::5.14:C;CHLE::HORSE::5.13:C;AMPC::ECOLI::5.05:C;SO1A1::RAT::5.03:C;MDR1B::MOUSE::5.:C;ADA1D:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;KCNK6:::inh::D;KCNK1:::inh::D|CP2D6:::inh:8.7:DC;CP2C8:::inh::D;CP2C9:::inh::D;CP2B6:::inh::D;CP1A1:::inh::D;CP2E1:::sub::D;CP1A2:::inh::D;CP3A7:::sub::D;CP3A4:::inh::D|MDR1:::inh:6.37:DC;ABCBB:::inh::D;SO1B1:::inh::D;S22A4:::inh::D;MRP2:::inh::D;S22A8:::inh::D;SO1A2:::inh::D;S22A5:::inh::D;S22A1:::inh::D;S22A2:::inh::D|A1AG1
Zonisamide|ok_inv|CAH9:::inh:8.3:DC;CAH2:::inh:7.99:DC;CAH5A:::inh:7.7:DC;CAH5B:::inh:7.69:DC;CAN::CANAL::7.46:C;CAH1:::inh:7.25:DC;CAH6:::inh:7.05:DC;CAN::YEAST::6.97:C;CAH7:::inh:6.93:DC;CYNT::HELPY::6.66:C;CAH13:::inh:6.37:DC;CAH15::MOUSE::6.2:C;MTCA2::MYCTU::6.06:C;LMNA::::6.05:C;AOFB::RAT::5.54:C;AOFB:::inh:5.51:DC;CAH14:::inh:5.28:DC;CAH4:::inh:5.07:DC;CAH3::BOVIN::5.07:C;AOFA:::inh::D;CAH12:::inh::D;CAH11:::inh::D;CAH10:::inh::D;CAH8:::inh::D;CAH3:::inh::D;CAC1I:::inh::D;CAC1H:::inh::D;CAC1G:::inh::D;SCN4B:::inh::D;SCN3B:::inh::D;SCN2B:::inh::D;SCN1B:::inh::D;SCNBA:::inh::D;SCN9A:::inh::D;SCN5A:::inh::D;SCN4A:::inh::D;SCN3A:::inh::D;SCN2A:::inh::D;SCN1A:::inh::D|CP3A5:::sub::D;UD11:::sub::D;CP2CJ:::inh::D;AOXA:::sub::D;CP3A4:::sub::D||
Paricalcitol|ok_inv|VDR:::ago::D|UD14:::sub::D;CP3A4:::sub::D;CP24A:::sub::D||
Tinidazole|ok_inv|LMNA::::5.7:C;DNA:::bin::D|CP3A4:::sub::D|ABCBB:::sub::D|
Repaglinide|ok_inv|ABCC8:::inh:7.3:DC;LMNA::::6.4:C;MK01::::5.2:C;S22A1::::5.04:C;PPARG:::ago::D|CP2C8:::sub::D;CP3A4:::sub::D|ABCBB:::sub::D;SO1B1:::sub::D|ALBU
Anileridine|ok_ill|OPRM:::ago::D|||
Phenformin|ok_out|LMNA::::6.4:C;HIF1A::::5.2:C;TSHR::::5.1:C;KCNJ8:::inh::D;AAPK1:::act::D|CP2D6:::sub:5.:DC|S22A1:::sub:5.:DC;S22A2:::inh::D|
Amantadine|ok|SGMR1::::7.69:C;M2::I000F::6.49:C;NFKB1::::5.55:C;TSHR::::5.2:C;NMDZ1::::5.:C;ACHA3:::ant::D;ACHA4:::ant::D;DRD2:::ago::D;ACHA7:::ant::D;NMD3A:::ant::D;M2::I60A0:inh::D|AOFB:::inh::D;DDC:::ind::D|S22A1:::inh::D;S22A2:::inh::D|
Metronidazole|ok|LMNA::::5.6:C;THB::::5.15:C;AL1A1::::5.1:C;MK01::::5.05:C;Protozoal_DNA::UNK:inh::D;Anaerobic_bacterial_DNA::UNK:inh::D;RDXA::HELPY:pot::D|CP3A7:::sub::D;CP3A5:::sub::D;CP2A6:::sub::D;UD11:::sub::D;CP2C8:::inh::D;CP3A4:::inh::D;CP2C9:::inh::D|MDR1:::inh::D|
Dinoprostone|ok|PE2R4:::ago:9.77:DC;PE2R2::RAT::9.7:C;PE2R3:::ago:9.48:DC;PE2R4::RAT::9.15:C;PE2R1:::ago:8.96:DC;PE2R2:::ago:8.77:DC;PE2R4::MOUSE::8.51:C;PE2R3::MOUSE::8.3:C;PE2R1::MOUSE::8.22:C;TSHR::::8.:C;PE2R2::MOUSE::7.66:C;MK01::::7.:C;PF2R::::6.6:C;PI2R::::6.59:C;S22A6::MOUSE::5.47:C;PD2R2:::ago::D||SO1B1:::sub::D;SO3A1:::sub::D;SO1C1:::sub::D;SO4A1:::sub::D;SO2A1:::sub::D;OSTB:::sub::D;OSTA:::sub::D;SO1A2:::sub::D;SO2B1:::sub::D;MRP4:::sub::D;S22A7:::inh::D;S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D;MRP5:::inh::D;S22A2:::inh::D|
Almotriptan|ok_inv|LMNA::::5.35:C;5HT1D:::ago::D;5HT1B:::ago::D|CP2C8:::sub::D;CP2E1:::sub::D;CP2CJ:::sub::D;FMO3:::sub::D;AOFA:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D||
Spectinomycin|ok_inv_vet|RS12::ECOLI:inh::D|||
Ketotifen|ok|HRH1:::ant:9.86:DC;HRH1::CAVPO::9.51:C;LMNA::::8.7:C;5HT2A::::8.05:C;5HT2B::::7.54:C;5HT2C::::7.08:C;ACM4::::6.85:C;ACM1::RAT::6.75:C;ACM1::::6.57:C;ACM5::::6.57:C;ACM2::::6.53:C;ADA2B::::6.49:C;LEF::BACAN::6.4:C;DRD1::::6.36:C;ACM3::::6.33:C;5HT6R::::6.28:C;DRD3::::6.18:C;ADA2A::::6.09:C;5HT1A::RAT::5.84:C;CP3A4::::5.8:C;ADA1D::::5.74:C;CP2D6::::5.5:C;TSHR::::5.4:C;HRH2::::5.39:C;6PGD:::inh::D|||
Buprenorphine|ok_ill_inv_vet|OPRM:::pag:8.8:DC;OPRM::MOUSE::8.44:C;OPRX;OPRD:::ant::D;OPRK:::ant::D|CP2CJ:::inh::D;CP2CI:::sub::D;CP2D6:::inh::D;CP3A7:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D;CP3A5:::sub::D;CP3A4:::inh::D|ABCG2:::inh::D;MDR1:::inh::D|
Levosimendan|ok_inv|PDE3A:::inh:8.1:DC;KCNJ8:::ind::D;KCJ11:::ind::D;TNNC1:::pot::D|||
Ceforanide|ok|Penicillin_binding_protein_2::BACFG:inh::D|||
Cyclobenzaprine|ok|ACM1::RAT::7.5:C;RET::::6.52:C;TSHR::::5.1:C;AOXA:::inh::D;TLR4:::inh::D;5HT7R:::ant::D;SC6A2:::inh::D;SC6A4:::inh::D;5HT6R:::ant::D;5HT2C:::ant::D;5HT2B:::ant::D;5HT2A:::ant::D|CP2D6:::sub:5.4:DC;UDB10:::sub::D;UD14:::sub::D;CP1A2:::sub::D;CP3A4:::sub::D||ALBU:::sub::D
Phenoxybenzamine|ok|ADA1B::RAT::8.74:C;DRD5::RAT::6.92:C;ADA1D:::ant::D;ADA1B:::ant::D;ADRB2;CALM1:::inh::D;ADA2B:::ant::D;ADA2C:::ant::D;ADA2A:::ant::D;ADA1A:::ant::D||S22A1:::inh:5.57:DC;S22A2:::inh:5.31:DC;S22A3:::inh:5.21:DC|
Etretinate|out|RARG:::ago::D;RXRB:::ago::D;RXRG:::ago::D;RARB:::ago::D;RXRA:::ago::D;RARA:::ago::D|CP19A:::inh::D||RABP1
Famotidine|ok|BLM::::8.8:C;HRH2::CAVPO::7.74:C;LMNA::::7.55:C;HRH2:::ant:7.39:DC;S47A1::::6.12:C;CYSP::TRYCR::5.:C||S22A8:::inh::D;S22A2:::inh::D|
Azacitidine|ok_inv|BLM::::8.8:C;MTOR::::6.93:C;ACM1::RAT::5.95:C;HBB::::5.9:C;LMNA::::5.8:C;NFKB1::::5.65:C;GEMI::::5.5:C;P53::::5.5:C;TPO::::5.5:C;AMPC::ECOLI::5.:C;DNA;RNA;DNMT1:::inh::D|CDD:::sub::D||
Misoprostol|ok|LMNA::::6.1:C;PE2R1:::ago::D;PE2R4:::ago::D;PE2R2:::ago::D;PE2R3:::ago::D|||
Colesevelam|ok|Bile_acids:::bin::D|||
Metacycline|ok_inv|MDFA::ECOLI::5.6:C;16S_ribosomal_RNA::Gut_flora:inh::D|||ALBU
Tipranavir|ok_inv|FACE1::MOUSE::5.92:C;PEPA5::::5.7:C;CATE::::5.05:C;Pol_polyprotein::9HIV1:inh::D|UD11:::ind::D;CP2CJ:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D|SO1B3:::inh::D;SO1B1:::inh::D;SO2B1:::inh::D;ABCBB:::inh::D|
Mesoridazine|ok_inv|KCNH2::::6.5:C;DRD2:::ant::D;5HT2A:::ant::D|CP2D6:::sub::D||
Maprotiline|ok_inv|HRH1:::ant:8.99:DC;SC6A2:::inh:7.92:DC;5HT2A:::bin:7.74:DC;5HT2C:::bin:7.39:DC;ACM4:::ant:7.24:DC;ADA1B::RAT::7.05:C;ACM3:::ant:7.:DC;ACM5:::ant:6.94:DC;ADA2B::::6.88:C;ACM1:::ant:6.84:DC;DRD1::::6.73:C;ADA1D::::6.71:C;5HT2B::::6.67:C;DRD3::::6.66:C;ADA1A::RAT::6.64:C;HRH2::::6.41:C;5HT6R::::6.38:C;DRD5::::6.37:C;ADA2C::::6.35:C;MTOR::::6.28:C;DRD2:::bin:6.18:DC;ADA2A,ADA2B,ADA2C:::ant:6.16,6.88,6.35:DC;ADA2A::::6.16:C;ACM2:::ant:6.16:DC;ACM1::RAT::5.65:C;SC6A3::::5.64:C;CP3A4::::5.6:C;LEF::BACAN::5.3:C;IMPA1::RAT::5.1:C;RORG::MOUSE::5.:C;5HT7R:::ant::D;ADA1A,ADA1B,ADA1D:::ant:,,6.71:DC|CP2D6:::sub:5.4:DC;CP1A2:::sub::D||A1AG1
Oxymetazoline|ok_inv|ADA2A:::ago:9.54:DC;5HT1B::::9.52:C;5HT1D::::9.4:C;5HT1B::RAT::9.04:C;ADA2C:::ago:9.:DC;ADA2A::BOVIN::8.82:C;ADA2C::RAT::8.72:C;ADA1B::RAT::8.72:C;5HT1A::RAT::8.49:C;NISCH::::8.21:C;ADA1A::RAT::8.19:C;ADA1A::BOVIN::7.88:C;ADA1A:::ago:7.8:DC;ADA2A::PIG::7.68:C;ADA2B::MOUSE::7.48:C;CP2D6::::7.4:C;ADA1B::MESAU::6.69:C;5HT2C::::6.52:C;ADA1D::RAT::6.48:C;5HT2A::::6.44:C;LMNA::::6.4:C;ACM4::::6.34:C;ADA2B:::bin:6.24:DC;5HT6R::::6.11:C;ADA1B:::ago:6.08:DC;ACM5::::6.02:C;ADA1D:::ago:5.87:DC;5HT2B::::5.71:C;ACM1::RAT::5.25:C|||
Salicylic_acid|ok_inv_vet|CAH2::::5.15:C;CAH15::MOUSE::5.14:C;CAH12::::5.06:C;CAH1::::5.:C;AK1C1:::inh::D;PGH2:::inh::D;PGH1:::inh::D|CP2C9:::sub::D|S22A7:::sub::D;MOT1:::sub::D;SO2B1:::sub::D;S22AB:::inh::D;S22A8:::inh::D;S22AA:::inh::D;S22A6:::inh::D|ALBU
Diethylpropion|ok_ill|SC6A2:::inh::D;SC6A3:::inh::D|||
Salmeterol|ok|ADRB2:::ago:10.15:DC;ADRB2::CAVPO::8.57:C;ADRB1:::ago:6.6:DC;ADRB3:::ago:6.:DC;DRD3::::5.98:C|CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D||
Meclofenamic_acid|ok_vet|PGH2:::inh:7.96:DC;PGH1::SHEEP::7.3:C;PGH2::RAT::7.:C;PGH2::MOUSE::6.7:C;PGH1:::inh:6.69:DC;FABPL::RAT::6.59:C;TTHY::::6.32:C;AK1C3::::6.27:C;MK01::::5.5:C;AK1C1::::5.5:C;AK1C2::::5.06:C;FABPI::::5.05:C;KCNQ3;KCNQ2;LOX5:::inh::D||SO1C1:::inh::D;S22A6:::inh::D|THBG:::sub::D
Methantheline|ok_inv|CP2D6::::5.4:C;LMNA::::5.4:C;CP1A2::::5.:C;HRH2:::ant::D;ACM1:::ant::D|||
Hexafluronium|ok|CHLE:::inh::D|||
Cycrimine|ok|ACM1:::ant::D|||
Zalcitabine|ok_inv|CXCR4::::7.06:C;LMNA::::7.:C;TAU::::6.9:C;NFKB1::::6.1:C;Reverse_transcriptase_RNaseH::9HIV1:inh::D|DCK:::sub::D|S29A2;S29A1;S22A7:::sub::D;S22A6:::sub::D|ALBU
Demecarium|ok|ACES:::inh::D;CHLE:::inh::D|||
Acetylsalicylic_acid|ok_vet|BLM::::8.55:C;TSHR::::7.3:C;PGH1::SHEEP::6.52:C;PGH1::BOVIN::6.46:C;ACM1::RAT::5.65:C;PGH2:::inh:5.62:DC;PGH2::SHEEP::5.62:C;PGH1:::inh:5.38:DC;ITB3::::5.3:C;Cyclin_A::UNK:rdw::D;PCNA:::rdw::D;MYC:::rdw::D;CCND1:::rdw::D;MK01,MK15,MK03,MK04,MK06,MK07;IKKB;CASP3:::idw::D;CASP1:::idw::D;TSG6:::idw::D;IKBA:::inh::D;KS6A3:::inh::D;BIP:::bin::D;P53:::ace::D;EDNRA:::inh::D;AAPK1,AAPK2,AAKB1,AAKB2,AAKG1,AAKG2,AAKG3:::act::D;AK1C1:::inh::D|ARY2:::sub::D;UD16:::sub::D;CP2C9:::sub::D;CP2CJ:::ind::D|S22A8:::inh::D;MDR1:::sub_ind::D;S22A6:::inh::D|
Phenprocoumon|ok_inv|VKOR1:::inh::D|CP2C8:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D||ALBU;A1AG1
Fulvestrant|ok_inv|ESR1:::ant::D|UD11:::sub::D;CP3A4:::sub::D||
Mezlocillin|ok_inv|PBPA::CLOPE:inh::D;PBP3::STREE:inh::D;MRDA::ECOLI:inh::D|||
Felbamate|ok|KPYM::::8.:C;SMN::::7.4:C;ACM1::RAT::6.5:C;CP2D6::::6.1:C;NPSR1::::6.1:C;NMDE1:::ant::D;NMD3A:::ant::D;NMDE2:::ant::D|CP2C9:::inh::D;CP2E1:::sub::D;CP2CJ:::inh::D;CP3A4:::sub_ind::D||
Fexofenadine|ok_inv|BLM::::8.05:C;HRH1:::ant:7.82:DC;LMNA::::6.8:C||S22A8:::sub::D;MRP3:::sub::D;MRP2:::sub::D;SO1A2:::sub::D;SO2B1:::sub::D;SO1B3:::sub::D;SO1B1:::sub::D;MDR1:::sub::D|A1AG1,A1AG2:::sub::D;ALBU:::sub::D
Isoniazid|ok_inv|DYR::MYCTU::9.:DC;CP3A4::::5.4:DC;PERM::::5.33:C;LUCI::PHOPY::5.3:C;INHA::MYCTU:cov::D;KATG::MYCTU:::D|CP1A2:::inh:5.2:DC;CP2CJ:::inh:5.:DC;CP2A6:::inh::D;NAT::MYCTU:inh::D;ARY2:::sub::D;CP2D6:::inh::D;CP2C9:::inh::D;CP2E1:::duo::D;CP2C8:::inh::DC||ALBU
Naratriptan|ok_inv|5HT1D:::ago:8.8:DC;5HT1B:::ago:8.48:DC;5HT1A:::ago:7.35:DC;5HT1F:::ago::D|AOFA:::sub::D||
Rizatriptan|ok|5HT1D:::ago:8.52:DC;5HT1B:::ago:8.:DC;5HT1D::PIG::7.3:C;5HT1A::::6.85:C;5HT3A::RAT::5.4:C;5HT2A::RAT::5.2:C;5HT2C::::5.1:C;5HT2A::::5.1:C;5HT1F:::ago::D|AOFA:::sub::D||
Dirithromycin|exp|23S_ribosomal_RNA::Gut_flora:inh::D|CP3A4:::inh::D||
Netilmicin|ok_inv|16S_ribosomal_RNA::Gut_flora:inh::D;RS12::ECOLI:inh::D|||
Hydrocodone|ok_ill_inv|OPRM:::ago:8.02:DC;OPRK::::6.59:C;LMNA::::5.05:C;SGMR1:::lig::D;OPRD:::ago::D|CP2CJ:::sub::D;CP2B6:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D||
Norgestimate|ok_inv|RORG::MOUSE::5.3:C;ANDR:::pag::D;ESR1:::ago::D;PRGR:::ago::D|CP3A4:::sub_ind::D|MRP2:::sub::D|
Carboplatin|ok|DNA:::cov::D|XDH:::ind::D;PERM:::sub::D;GSTT1:::sub::D;MT1A:::sub::D;MT2:::sub::D;SODC:::inh::D;GSTP1:::sub::D;GSTM1:::sub::D;NQO1:::sub::D|COPT1:::sub::D;COPT2:::sub::D;ATP7A:::sub::D;ATP7B:::sub::D;ABCG2:::sub::D;MRP2:::sub::D|
Methylprednisolone|ok_vet|GCR:::ago:8.3:DC;HIF1A::::7.3:C;NR1I2::RAT::5.4:C;ANXA1:::ago::D|CP2C9:::ind::D;CP2CJ:::ind::D;CP2C8:::ind::D;CP2B6:::ind::D;CP1B1:::ind::D;CP2A6:::ind::D;CP3A4,CP343,CP3A5,CP3A7:::sub_ind::D;CP3A4:::sub_ind::D;DHI1,DHI2;AK1C1,AK1C2,AK1C3,AK1C4:::sub::D|MDR1:::sub_ind::D|ALBU:::bin::D
Pindolol|ok_inv|ADRB2:::pag:9.42:DC;ADRB1:::pag:9.28:DC;5HT1A::RAT::7.7:C;5HT1A:::ant:7.65:DC;ACM1::RAT::7.5:C;ADRB3:::ago:7.18:DC;5HT1B::RAT::7.1:C;LMNA::::6.9:C;CP3A4::::6.5:C;5HT1B::::5.59:DC;NFKB1::::5.3:C;AGAL::::5.:C|CP2D6:::inh::D||
Mepivacaine|ok_vet|SCNAA:::inh::D|||
Zaleplon|ok_ill_inv|GBRA1:::pot:6.54:DC;GBRG2::::5.79:C;TSPO|AOXA:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D||
Bromfenac|ok|PGH1:::inh:8.07:DC|PGH2:::inh:8.32:DC||
Apraclonidine|ok|ADA2A:::ago:8.72:DC;ADA2B::RAT::8.32:C;ADA2C::::7.52:C;ADA1A:::ago:6.74:DC;HCD2::::5.9:C;ADA2B:::ago::D|||
Ethiodized_oil|ok_inv||||
Telmisartan|ok_inv|AGTRA::RAT::9.64:C;AGTR2::::9.48:C;AGTR1:::ant:9.31:DC;AGTRB::RAT::8.52:C;CP2J2::::7.:C;PPARG:::pag:6.15:DC;SO1B3::::6.02:C;SO1B1::::5.99:C;NPSR1::::5.9:C;GLRA1::::5.49:C;PPARG::MOUSE::5.39:C;CP2C9::::5.32:C;ACE::::5.22:C|UD13:::sub::D;CP2CJ:::inh::D|ABCBB:::sub::D;ABCG2:::inh::D;MRP2:::inh::D;MDR1:::inh::D|
Desloratadine|ok_inv|HRH1:::ant:9.01:DC;5HT2A::::8.02:C;5HT2C::::7.8:C;5HT2B::::7.55:C;ACM2::::7.42:C;ACM4::::7.33:C;ACM1::::7.19:C;ACM3::::7.02:C;SC6A4::::6.91:C;ACM5::::6.68:C;GLRA2::RAT::6.33:C;DRD3::::6.19:C;ADA2B::::6.01:C;5HT6R::::6.:C;HRH2::::5.97:C;SC6A2::::5.96:C;ADA1B::RAT::5.7:C;SC6A3::::5.51:C;LMNA::::5.5:C||MDR1:::inh::D|
Methyldopa|ok|HCD2::::6.9:C;TYDP1::::6.3:C;KPYK::LEIME::6.1:C;DPOLB::::5.95:C;LOX15::::5.9:C;RECQ1::::5.85:C;LOX15::RABIT::5.67:C;KDM4E::::5.52:C;TAU::::5.5:C;BLM::::5.45:C;LYAG::::5.45:C;FYN::::5.29:C;EGFR::::5.28:C;AL1A1::::5.25:C;APEX1::::5.1:C;DDC:::inh::D;ADA2A|COMT:::sub::D|S15A1:::inh::D|
Alosetron|ok_out|5HT3A:::ant:9.3:DC;5HT2B::::7.19:C;KCNH2::::5.64:C|CP3A4:::sub:6.22:DC;CP1A2:::inh:6.22:DC;CP2E1:::inh::D;CP2C9:::sub::D||
Dactinomycin|ok_inv|RORG::MOUSE::7.75:C;HD::::7.5:C;HIF1A::::6.6:C;RECQ1::::5.85:C;CYSP::TRYCR::5.4:C;GRB2::::5.3:C;GRB2::MOUSE::5.3:C;BLM::::5.15:C;DDR2::::5.05:C;TOP2A,TOP2B:::inh::D;DNA:::cov::D||ABCG2:::sub::D;MRP1:::sub::D;MRP6:::sub::D;MDR1:::inh::D;S22A5:::inh::D|
Selenium_Sulfide|ok||||
Azelastine|ok|HRH1:::ant:9.7:DC;ADA1A::::7.3:C;ADA1B::::7.3:C;KCNH2::::7.:C;HRH3::::6.83:C;CAC1C::CAVPO::5.1:C;LTC4S:::inh::D;PA21B:::inh::D;HRH2:::inh::D|CP2D6:::inh:6.:DC;CP2B6:::inh::D;CP2E1:::inh::D;CP2A6:::inh::D;CP2C8:::sub::D;CP2C9:::inh::D;CP3A5:::sub::D;CP1A1:::inh::D;CP2CJ:::inh::D;CP1A2:::sub::D;CP3A4:::inh::D|MDR1:::inh::D|
Ezetimibe|ok|NPCL1::RAT::6.7:C;NPSR1::::5.3:C;RORG::MOUSE::5.15:C;AMPN;NPCL1:::inh::D;SOAT1:::inh::D|CP2C8:::inh::D;CP3A4:::inh::D;UD2B7:::sub::D;UDB15:::sub::D;UD13:::sub::D;UD11:::sub::D|ABCBB:::sub::D;ABCG8:::sub::D;ABCG2:::sub::D;MRP3:::sub::D;ABCG5:::sub::D;SO1B1:::sub::D;MRP2:::sub::D;MDR1:::sub::D|
Edetic_acid|ok_vet|Manganese_cation:::chel::D;Iron:::chel::D;Lead:::chel::D|CP19A:::sub::D;PON3:::inh::D;ADA:::inh::D||
Dipyridamole|ok|LMNA::::8.4:C;S29A1::::8.09:C;CNCG::::6.9:C;PDE11::::6.4:C;PDE4A:::inh:6.3:DC;PDE5A:::inh:6.28:DC;PDE7A::::6.22:C;PRUN1::::6.11:C;PDE10:::inh:6.:DC;CP2CJ::::5.9:C;TAU::::5.85:C;RORG::MOUSE::5.85:C;S22A2::::5.59:C;MEN1::::5.5:C;PDE2A::::5.49:C;CASP7::::5.4:C;CASP1::::5.4:C;NF2L2::::5.39:C;CP2C9::::5.3:C;NPSR1::::5.2:C;LOX15::RABIT::5.16:C;TPO::::5.:C;CP3A4::::5.:C;CP2D6::::5.:C;GNAI1::::5.:C;KMT2A::::5.:C;LEF::BACAN::5.:C;A1AG1;RCAN1;ADA:::inh::D||MRP4:::inh:5.7:DC;ABCBB:::sub::D;SO2B1:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;MDR1:::inh::D;MRP5:::inh::D|
Telithromycin|ok|23S_ribosomal_RNA::Gut_flora:inh::D|CP3A4:::inh::D|SO1B1:::inh:5.46:DC;SO1B3:::inh:5.23:DC|
Ethinylestradiol|ok|ESR1:::ago:9.89:DC;ST1A1::::8.37:C;ESR2::::8.09:C;SC6A4::::7.54:C;SHBG::::6.81:DC;AOXA::::6.37:C;SC6A3::::6.35:C;GCR::::6.11:C;CP2B6::::6.1:C;SC6A2::::6.02:C;ANDR::RAT::5.96:C;5HT4R::CAVPO::5.88:C;S22A2::::5.66:C;NR1I3::::5.52:C;LOX15::RABIT::5.25:C;NR1I2:::ago::D|CP2CJ:::inh::D;UD11:::sub_ind::D;CP2C8:::inh::D;CP3A4:::sub::D|MDR1:::sub::D;MRP2:::ind::D;NTCP:::ind::D;ABCBB:::duo::D|
Lomefloxacin|ok_inv|TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A2:::inh::D|MRP2:::inh::D;S22A5:::inh::D|
Cyclopentolate|ok|ACM1:::ant::D|CHLE:::sub::D||
Ramelteon|ok_inv|MTR1A::::10.86:DC;MTR1B::::10.35:DC|CP2C9:::sub::D;CP3A4:::sub::D;CP2CJ:::sub::D;CP1A2:::sub::D||
Physostigmine|ok_inv|ACES:::inh:9.37:DC;ACES::MOUSE::9.17:C;ACES::RAT::9.17:C;ACES::ELEEL::9.:C;LMNA::::8.4:C;ACES::TETCF::7.96:C;CHLE::HORSE::7.85:C;CHLE::::7.82:C;ACES::CHICK::7.7:C;ACES::BOVIN::7.52:C;CP2D6::::6.7:C;BLM::::6.55:C;CHLE::MOUSE::6.55:C;ACHB2;ACHA4|||
Isotretinoin|ok|MK01::::6.34:C;5HT2B::::6.27:C;RABP1::CHICK::6.05:C;AA3R::::5.63:C;PMP22::::5.62:C;MK14::::5.6:C;ADA2B::::5.52:C;MTOR::::5.33:C;RARG;RARA|CP3A4:::sub::D||ALBU:::bin::D
Formoterol|ok_inv|ADRB2:::ago:9.72:DC;ADRB2::CAVPO::9.4:C;ADRB1:::ago:7.9:DC;ADRB3:::ago:7.6:DC;DRD3::::5.79:C|CP2A6:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP2D6:::sub::D||
Nandrolone_phenpropionate|ok_ill_inv|ANDR:::ago::D|||
Dimenhydrinate|ok|LMNA::::9.:C;HRH1:::ant:7.43:DC;ACM4::::7.1:C;ACM3::::7.02:C;ACM1::::6.96:C;ACM2::::6.79:C;5HT2A::::6.7:C;ACM5::::6.64:C;5HT2C::::6.48:C;SGMR1::::6.31:C;5HT2B::::5.96:C;ADA1D::::5.85:C;CP2D6::::5.82:C;ADA2A::::5.79:C;SC6A3::::5.75:C;SC6A2::::5.69:C;ADA2B::::5.6:C;CP1A2::::5.3:C|||
Glycopyrronium|ok_inv_vet|ACM1:::ant:9.9:DC;ACM4::::9.8:C;ACM5::::9.7:C;ACM3:::ant:9.6:DC;ACM2:::bin:9.3:DC|||
Cytarabine|ok_inv|LMNA::::7.4:C;MTOR::::7.13:C;LMP1::EBVB9::6.13:C;NCOA3::::5.12:C;DNA:::cov::D;DPOLB:::inh::D|DCTD:::sub::D;5NTD:::sub::D;DCK:::sub::D;CP3A4:::sub::D;CDD:::sub::D|S29A1:::sub::D;MRP7:::sub::D;S22A4:::sub::D|
Dopamine|ok|DRD2:::ago:9.16:DC;DRD2::RAT::8.96:C;DRD4:::ago:8.92:DC;DRD3:::ago:8.74:DC;DRD2::BOVIN::8.74:C;DRD5::RAT::8.7:C;DRD4::RAT::8.62:C;DRD1::BOVIN::8.43:C;SC6A2:::inh:8.18:DC;DRD3::RAT::7.96:C;DRD1,DRD5:::ago:7.7,5.61:DC;DRD1:::ago:7.7:DC;ADA2C::RAT::7.24:C;DRD1::RAT::6.82:C;SC6A3::RAT::6.7:C;TYDP1::::6.35:C;SC6A3:::ind:6.34:DC;HCD2::::6.3:C;AA2BR::RAT::6.01:C;FFP::BACIU::5.9:C;TAU::::5.8:C;RECQ1::::5.75:C;DRD5:::ago:5.61:DC;ADA1A::::5.6:C;KDM4E::::5.52:C;SGMR1::RAT::5.52:C;TPO::::5.5:C;ARP19::RAT::5.46:C;MTR1A::::5.15:C;MTR1B::::5.04:C;ADRB1::RAT::5.:C;HIF1A::::5.:C;VMAT2;SODC;5HT3B;5HT3A;SC6A4:::inh::D;5HT7R:::bin::D;5HT1A:::bin::D|COMT:::sub::D;AOFB:::sub::D;AOFA:::sub::D;DOPO:::sub::DC|PO5F1:::sub::D;S22A5:::inh::D;S22A3:::inh::D;S22A1:::sub::D;S22A2:::inh::D|
Rivastigmine|ok_inv|CHLE:::inh:7.52:DC;ACES:::inh:7.43:DC;ACES::BOVIN::6.21:C;CHLE::HORSE::6.08:C;ACES::MOUSE::5.95:C;CHLE::MOUSE::5.8:C;ACES::RAT::5.74:C;ACES::ELEEL::5.47:C|||
Exemestane|ok_inv||CP19A:::inh:7.99:DC;CP3A4:::sub::D||
Oxaprozin|ok|LMNA::::6.45:C;PGH1:::inh:6.07:DC;LEF::BACAN::5.3:C;MK01::::5.3:C;PGH2:::inh::D|||
Methyl_aminolevulinate|ok_inv|FCGR1:::abo::D|||
Azathioprine|ok|BLM::::6.7:C;HBB::::6.5:C;LMNA::::6.4:C;P53::::6.1:C;GEMI::::5.75:C;CP3A4::::5.4:C;ACM1::RAT::5.:C;RAC1;HPRT:::inh::D|CP1A2:::sub::D;GSTM1:::sub::D;GSTA2:::sub::D;GSTA1:::sub::D;TPMT:::sub::D;XDH:::sub::D||
Neomycin|ok_vet|RS12::ECOLI:inh::D;16S_ribosomal_RNA::Gut_flora:inh::D;CASR|||
Auranofin|ok_inv|PRDX5:::inh::D;IKKB:::inh::D|||ALBU
Gabapentin|ok_inv|CA2D1:::inh:7.57:DC;CA2D1::MOUSE::6.92:C;CA2D1::RAT::5.05:C;KCNQ5:::act::D;KCNQ3:::act::D;AA1R:::ago::D;A0A024R8I1,CAC1B::,HUMAN:inh::D;CA2D2:::inh::D|BCAT1:::inh::D|LAT1:::sub::D|
Doxorubicin|ok_inv|AURKA::::7.4:C;HIF1A::::6.92:C;EBP::::6.82:C;TOP2A:::inh:6.:DC;MMP2::::5.96:C;5HT4R::CAVPO::5.68:C;ERBB2::::5.6:C;CISD1::::5.46:C;ACM1::::5.43:C;FYN::::5.29:C;NOLC1;DNA:::itc::D|NCPR:::sub::D;NDUS7:::sub::D;NDUS3:::sub::D;NDUS2:::sub::D;NOS3:::sub::D;NOS2:::sub::D;NOS1:::sub::D;XDH:::sub::D;NQO1:::sub::D;AK1C3:::sub::D;AK1A1:::sub::D;CBR3:::sub::D;CBR1:::sub::D;CP1B1:::duo::D;CP2B6:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D|MDR1:::duo:5.07:DC;MRP2:::sub::D;RBP1:::sub::D;ABCBB:::sub::D;ABCB8:::sub::D;MRP7:::inh::D;S22AG:::sub::D;ABCG2:::sub::D;MRP6:::inh::D;MRP3:::inh::D;MRP1:::inh::D|ALBU
Frovatriptan|ok_inv|5HT1D:::ago:8.36:DC;5HT1B:::ago:7.99:DC;5HT1A::::7.21:C|CP1A2:::sub::D||
Hydrochlorothiazide|ok_vet|LMNA::::8.35:C;THB::::6.55:C;CAH2::::6.54:C;CAH1::::6.48:C;KCMA1:::inh::D;S12A3:::inh::D||MRP4:::sub::D;S22AB:::sub::D;S22A8:::sub::D;S22A6:::inh::D|ALBU:::bin::D
Cyclacillin|ok|LMNA::::5.9:C;PBP2A::STAAU:inh::D;PBP3::STREE:inh::D;PBPA::STRR6:inh::D;PBPA::CLOPE:inh::D||S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|
Salbutamol|ok_vet|ADRB2::CAVPO::9.34:C;ADRB2:::ago:7.6:DC;ADRB2::BOVIN::6.28:C;ADRB3;ADRB1:::ago::D|CP3A4:::inh::D||
Levobupivacaine|ok_inv|IMPA1::RAT::8.:C;CP2D6::::6.71:C;TSHR::::5.2:C;SCNAA:::inh::D|CP1A2:::sub:5.3:DC;CP3A4:::sub:5.:DC||
Cromoglicic_acid|ok|GPR35::::6.68:C;LMNA::::6.15:C;TYDP1::::5.75:C;S100P:::ant::D;KCMA1:::inh::D|||
Ganciclovir|ok_inv|BLM::::8.49:C;LMNA::::5.5:C;HIF1A::::5.4:C;NFKB1::::5.:C;MEN1::::5.:C;KITH::HHV11:ind::D;DNA:::destbz::D;DPOL::HHV11:inh::D||S47A2:::sub::D;S47A1:::sub::D;S22A7:::inh::D;S22A8:::inh::D;S22A6:::inh::D;S22A1:::inh::D|
Hydroxyurea|ok|NFKB1::::5.5:C;RIR1:::inh::D|CP2D6:::inh::D||
Letrozole|ok_inv|C11B2::::5.85:C;C11B1::::5.58:C;CP2CJ::::5.1:C;TSHR::::5.1:C|CP19A:::inh:10.7:DC;CP3A4:::sub:5.3:DC;CP2A6:::inh::D||
Tioconazole|ok|CP17A::::6.3:C;CP51A:::inh::D;CP51::CANAL:ant::D|CP3A4:::inh::D;CP2E1:::inh::D;CP2CJ:::inh::D;CP19A:::inh::D||
Busulfan|ok_inv|LMNA::::6.1:C;MMP9::::5.28:C;DNA:::cov::D|MGST2:::sub::D;GSTP1:::sub::D;GSTM1:::sub::D;GSTA1:::sub::D;GSTA2:::sub::D;CP3A4:::sub::D||
Ketoprofen|ok_vet|PGH1:::inh:8.7:DC;PGH2:::inh:7.59:DC;SMN::::7.3:C;PGH1::SHEEP::7.17:C;LMNA::::6.5:C;S22A6::RAT::6.3:C;S22A7::RAT::5.74:C;AMPC::ECOLI::5.45:C;TAU::::5.4:C;MK01::::5.05:C;CXCR1|UD11:::sub::D;CP2C8:::inh::D;CP2C9:::inh::D|S22A6:::inh:5.89:DC;S22A7:::inh::D;S22AB:::inh::D;S22A8:::inh::D;SO1A2:::inh::D;MRP4:::inh::D|ALBU
Edrophonium|ok|CHLE:::inh::D;ACES:::inh::D|||
Metyrapone|ok_inv|C11B1::BOVIN::6.24:C;C11B1::RAT::5.34:C;LMNA::::5.1:C;CPXA::PSEPU:::D|C11B2:::inh:8.3:DC;C11B1:::inh:7.84:DC;CP3A4:::duo:6.1:DC;CP2E1:::inh::D;CP2A6:::inh::D|MRP3:::ind::D|
Cinacalcet|ok|CASR:::ago:7.1:DC;GLRA1::::6.49:C|CP2D6:::inh:7.3:DC;CP1A2:::sub::D;CP3A4:::sub::D||
Clobetasol_propionate|ok|GCR:::ago:9.18:DC;GCR::RAT::8.5:C;NPSR1::::6.:C;ANDR::RAT::5.6:C;ABCBB::::5.07:C|CP3A5:::ind::D;CP3A4:::sub_ind::D||
Balsalazide|ok_inv|LOX5:::inh::D;PGH1:::inh::D;PGH2:::inh::D;PPARG:::ago::D|AZRB::BACOY:sub::D||
Sulfamethoxazole|ok|DYR::PNECA::7.:C;EDNRA::RAT::5.4:C;DHPS::ECOLI:inh:5.33:DC;TAU::::5.05:C;GSTP1|CP3A4:::sub::D;CP2C8:::inh::D;UD19:::sub::D;PGH1:::sub::D;CP2C9:::inh::D;ARY2:::sub::D;ARY1:::sub::D|ABCBB:::sub::D|ALBU
Glyburide|ok|KCJ11,KCNJ8:::inh:8.37,:DC;KCJ11::::8.37:C;TSHR::::6.9:C;SO1B1::::5.85:C;S22A6::RAT::5.8:C;CISD1::::5.78:C;HIF1A::::5.7:C;ABCBB::RAT::5.55:C;S15A2::RAT::5.11:C;CP2D6::::5.:C;TRPM4:::inh::D;CFTR:::ant::D;CPT1A:::inh::D;ABCA1:::inh::D;ABCC9:::mod::D;ABCC8,KCJ11:::inh:,8.37:DC|CP2C9:::inh:5.8:DC;CP3A4:::inh:5.4:DC;CP2CJ:::sub:5.:DC;CP3A5:::sub::D;CP3A7:::sub::D|ABCBB:::inh:5.28:DC;SO2B1:::sub::D;S22A7:::inh::D;ABCG2:::sub::D;MRP2:::inh::D;S22A6:::inh::D;S15A2:::inh::D;SO1A2:::inh::D;S15A1:::inh::D;MRP1:::inh::D;MDR1:::inh::D;MRP3:::inh::D|ALBU:::bin::D
Minocycline|ok_inv|MDFA::ECOLI::5.59:C;CYC:::neg::D;CASP3:::neg::D;CASP1:::neg::D;VEGFA:::inh::D;MMP9:::inh::D;LOX5:::inh::D;IL1B:::mod::D;16S_ribosomal_RNA::Gut_flora:inh::D;RS4::ECOLI:inh::D;RS9::ECOLI:inh::D||S22A7:::inh::D;S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D|
Guanfacine|ok_inv|ACM1::RAT::7.9:C;NISCH::::7.72:C;ADA2A:::ago:7.3:DC;ADA2B:::bin:6.94:DC;CP2D6::::6.9:C;LMNA::::6.45:C;ADA1A::RAT::6.26:C;5HT2C::::6.12:C;5HT2A::::6.06:C;ADA2C::::6.03:C;5HT2B::::5.87:C;HCD2::::5.1:C;HIF1A::::5.:C|CP2CJ:::sub:6.6:DC;CP3A4:::sub::D||
Bethanechol|ok|ACM3::::7.01:DC;ACM4;ACM1;ACM2:::ago::D|||
Isosorbide_mononitrate|ok|GCYA2:::ind::D|||
Trichlormethiazide|ok_vet|CAH7::::8.1:C;CAH9::::7.06:C;CAH2:::inh:7.04:DC;CAH5B::::6.87:C;CAH12::::6.51:C;CAH1:::inh:6.46:DC;CAH4:::inh:6.35:DC;CAH13::MOUSE::6.19:C;CAH5A::::6.12:C;CAH6::::5.61:C;CAH14::::5.46:C;AT1A1:::inh::D;S12A3:::inh::D|TPMT:::inh::D||
Phylloquinone|ok_inv|OSTCN:::ago::D;VKGC:::ind::D|||
Felodipine|ok_inv|AA3R::::6.22:C;NR1I2::::5.72:C;NR1H4::::5.3:C;TNNC1;TNNC2;MCR:::ant::D;PDE1A:::inh::D;PDE1B:::inh::D;CALM1;CA2D2:::inh::D;CAC1H:::inh::D;CAC1S:::inh::D;CAC1D:::inh::D;CACB2:::inh::D;CA2D1:::inh::D;CAC1C:::inh::D|CP2C9:::inh:5.34:DC;CP2D6:::inh::D;CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::inh::D|ABCBB:::sub::D;MDR1:::inh::D|
Mycophenolic_acid|ok|IMDH2:::inh:8.22:DC;IMDH1:::inh:7.72:DC;SMN::::7.2:C;LMNA::::6.85:C;LEF::BACAN::5.9:C;KDM4E::::5.05:C;CP3A4::::5.:C|UD2B7:::sub:5.82:DC;UD16:::sub::D;UD17:::sub::D;UD19:::sub::D;UD11:::sub::D||
Amlexanox|ok_out|NPC1::::6.5:C;RAB9A::::6.3:C;RORG::MOUSE::5.4:C;KPYK::LEIME::5.15:C;FGF1:::inh::D;IL3:::ant::D;S10AD:::ant::D;S10AC:::ant::D|||
Ketoconazole|ok_inv|C11B2::::7.17:C;CP17A:::inh:7.09:DC;NR1I3;NR1I2:::ant::D;KCNH2:::inh::D;CP21A:::inh::D;ANDR:::bin::D;CP51::CANGA:inh::D|CP3A4:::inh:7.92:DC;CP3A5:::inh:6.92:DC;C11B1:::inh:6.9:DC;CP4F2:::inh::D;CP19A:::inh::D;CP4FC:::inh::D;UD2B7:::inh::D;UD17:::inh::D;UD11:::inh::D;CP2D6:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;CP2B6:::inh::D;CP1B1:::inh::D;CP2A6:::inh::D;CP1A2:::inh::D;CP1A1:::duo::D;CP2CJ:::inh::D|SO1B1:::inh::D;MDR1:::inh::D;ABCBB:::inh::D|SHBG:::lig::D;ALBU:::lig::D
Methoxyflurane|ok_inv_vet|GABAR:::aga::D;NU1M;ATPD;KCNA1:::ind::D;AT2C1:::inh::D;GLRA1:::ago::D;GRIA1:::ant::D;GBRA1:::ago::D|CP3A4:::sub::D;CP2D6:::sub::D;CP2C9:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;CP1A2:::sub::D;CP2E1:::sub::D||
Irbesartan|ok_inv|AGTR1:::ant:9.1:DC;AGTRB::RAT::9.1:C;LMNA::::6.4:C;LYAG::::6.35:C;EDNRA::::5.:C;JUN|CP3A4:::inh::D;PGH1:::sub::D;UD13:::sub::D;CP2C9:::sub::D;CP2C8:::inh::D||A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Topotecan|ok_inv|HIF1A::::7.92:C;TOP1:::inh:7.58:DC;DNA:::itc::D;TOP1M:::inh::D|CP3A4:::duo:5.82:DC|S47A1:::inh:5.89:DC;S47A2:::sub:5.07:DC;MDR1:::sub::D;ABCG2:::sub::D|
Ethinamate|ok_ill_out|CAH1:::inh::D;CAH2:::inh::D|||
Probenecid|ok_inv|CAH9::::6.44:C;CAH2::::6.37:C;CAH12::::5.9:C;S22A8::MOUSE::5.52:C;S22A8::RAT::5.35:C;S22A6::MOUSE::5.2:C;S22AK::MOUSE::5.08:C;T2R16;PANX1:::ant::D|CP2C9:::inh::D;UD11:::inh::D;CP3A4:::ind::D;CP2C8:::ind::D|S22A6:::inh:5.37:DC;S22A8:::inh:5.36:DC;GTR9:::inh::D;S22AC:::inh::D;S22A7:::inh::D;SO1C1:::inh::D;ABCCB:::inh::D;MRP2:::inh::D;S22AA:::inh::D;NTCP:::inh::D;MOT1:::inh::D;SO1A2:::inh::D;MRP1:::inh::D;MRP6:::inh::D;S22A5:::inh::D;MOT2:::inh::D;MRP5:::inh::D;MRP4:::inh::D;MRP3:::inh::D;S22A1:::inh::D;S22A2:::inh::D;S22AB:::inh::DC|ALBU
Mercaptopurine|ok|HBB::::5.5:C;AL1A1::::5.1:C;P53::::5.1:C;IMDH1,IMDH2:::inh::D;PUR1:::inh::D;HPRT:::inh::D|AOXA:::sub::D;XDH:::sub::D;TPMT:::sub::D|S29A2:::sub::D;S29A1:::sub::D;S28A3:::sub::D;S28A2:::sub::D;MRP5:::sub::D;MRP4:::sub::D;S22A8:::inh::D|
Procainamide|ok|LMNA::::8.:C;ACES::BOVIN::6.3:C;ACES::::6.:C;S22A1::MOUSE::5.41:C;ACM1::RAT::5.2:C;S22A1::RAT::5.15:C;KCNH2:::inh::D;DNMT1;SCN5A:::inh::D|CHLE:::inh::D;CP2D6:::sub::D|S47A2:::sub::D;S47A1:::sub::D;S22A4:::inh::D;S22A5:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|
Tolterodine|ok_inv|ACM1:::ant:8.85:DC;ACM5:::ant:8.66:DC;ACM2:::ant:8.57:DC;ACM4:::ant:8.51:DC;ACM3:::ant:8.49:DC;ACM2::RAT::8.16:C;ACM3::RAT::8.15:C;KCNH2::::7.9:C;CAC1C::CAVPO::6.84:C;TAU::::5.3:C;RORG::MOUSE::5.25:C;SCN5A::::5.2:C|CP2CJ:::sub::D;CP2C9:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D||
Selegiline|ok_inv_vet|AOFB:::inh:10.77:DC;AOFB::RAT::8.56:C;AOFA::RAT::7.74:C;AOFA:::inh:7.17:DC;ADA2B::::6.76:C;ADA2A::::6.17:C;AOFB::BOVIN::6.01:C;CP2B1::RAT::5.98:C;AOFA::BOVIN::5.42:C|CP2E1:::inh::D;CP2D6:::inh::D;CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1A2:::inh::D;CP2A6:::inh::D;CP3A4:::sub::D;CP2B6:::inh::D|MDR1:::inh::D|
Fenofibrate|ok|FABPL::RAT::7.74:C;ACM1::RAT::7.2:C;PPARG::::6.24:C;5HT2A::::6.22:C;PPARA:::ago:6.:DC;5HT2C::::5.91:C;AA3R::::5.49:C;TYDP1::::5.45:C;CP3A4::::5.4:C;TAU::::5.35:C;CP1A2::::5.3:C;UBP2::::5.2:C;SC6A3::::5.16:C;MEN1::::5.05:C;NR1I2:::pag::D;MMP25:::inh::D|CP2C9:::inh:5.3:DC;CP2CJ:::inh:5.1:DC;ALDR:::sub::D;AK1C3:::sub::D;AK1C2:::sub::D;AK1C1:::sub::D;CP2A6:::inh::D;CP2C8:::inh::D;CBR1:::sub::D;EST1:::sub::D;UD19:::sub::D|ABCBB:::sub::D|ALBU:::bin::D
Thalidomide|ok_out|PGH1::SHEEP::6.43:C;PGH2::SHEEP::6.3:C;A1AG1,A1AG2:::bin::D;FGFR2:::ant::D;DNA:::itc::D;NFKB1:::ant::D;TNFA:::inh::D;CRBN:::inh::D|CP3A5:::ind::D;PGH1:::sub::D;CP2C9:::sub::D;CP2E1:::sub::D;CP1A1:::sub::D;CP2CJ:::inh::D;PGH2:::sub::DC||
Melphalan|ok|AL1A1::::5.55:C;CP3A4::::5.5:C;FFP::BACIU::5.25:C;DNA:::cov::D||LAT1;S22A3:::inh::D|
Memantine|ok_inv|NMDZ1:::bin:9.02:DC;NMDE3::RAT::6.15:C;NMDZ1::RAT::5.96:C;MTOR::::5.18:C;GLRA1,GLRA2,GLRA3,GLRA4,GLRB:::inh::D;GABAR:::bin::D;NMDA:::ant::D;DRD2:::duo::D;Alpha_7_nicotinic_cholinergic_receptor_subunit:::ant::D;5HT3A:::ant::D|CP2CJ:::inh::D;CP2A6:::inh::D;CP2B6:::inh::D|S47A1;S22A4;SL9A1;S22A2:::sub::D|
Gatifloxacin|ok_inv|GYRB::ECOLI::6.3:C;STRP::STRP1::6.18:C;PARC::STAAU::5.92:C;CLK4::::5.4:C;CLK2::::5.1:C;KPCD3::::5.1:C;GYRA::MYCTU::5.03:C;PARE::STRPN:inh::D;PARC::STRPN:inh::D;GYRB::STRPN:inh::D;GYRA::STRPN:inh::D|CP1A2:::inh::D||ALBU
Rifampicin|ok|INHA::MYCTU::7.52:C;NR1I2:::ago:6.72:DC;SO1A4::RAT::5.85:C;LOX15::RABIT::5.53:C;CASP1::::5.08:C;RPOB::ECOLI:inh::D|CP2B6:::ind:5.89:DC;CP3A5:::ind::D;UD19:::inh::D;CP3A7:::ind::D;CP343:::ind::D;CP2E1:::ind::D;CP2A6:::ind::D;CP2CJ:::ind::D;UD11:::ind::D;CP3A4:::ind::D;CP2C8:::ind::D;CP1A2:::ind::D;CP2C9:::ind::D|SO1B1:::inh:6.52:DC;SO1B3:::inh:5.85:DC;S22A8:::inh::D;S22A6:::inh::D;MRP2:::ind::D;ABCBB:::inh::D;SO1A2:::inh::D;SO2B1:::inh::D;MRP5:::ind::D;MRP3:::ind::D;S22A7:::inh::D;MRP1:::inh::D;MDR1:::ind::D|A1AG1,A1AG2:::lig::D;ALBU:::lig::D
Lubiprostone|ok_inv|CLCN2:::ind::D|CBR1:::sub::D||
Fluocinonide|ok_inv|HIF1A::::9.:C;GCR:::ago:8.62:DC;SMO:::ago::D|CP3A5:::ind::D;CP3A4:::sub_ind::D||CBG:::bin::D
Abacavir|ok_inv|HLAB;Reverse_transcriptase_RNaseH::9HIV1:inh::D|ADK:::sub::D;UD11:::sub::D;ADH6:::sub::D||
Ergoloid_mesylate|ok|DRD1:::duo::D;ADA1A:::duo::D;ADRB1:::duo::D;5HT1A:::duo::D|CP3A4:::sub::D||
Ibuprofen|ok|LMNA::::8.25:C;PGH2:::inh:7.:DC;PGH1:::inh:6.67:DC;PGH1::MOUSE::6.66:C;NFKB1::::6.65:C;PGH2::MOUSE::6.07:C;PGH1::SHEEP::5.97:C;PGH2::SHEEP::5.96:C;S22AK::MOUSE::5.96:C;PGH2::BOVIN::5.96:C;ALBU::RAT::5.83:C;PGH2::RAT::5.7:C;PGH1::BOVIN::5.54:C;ALBU::BOVIN::5.52:C;S22A6::RAT::5.46:C;S22A6::MOUSE::5.33:C;S10A7:::ind::D;GP1BA:::ind::D;PPARA:::act::D;CFTR:::inh::D;PPARG:::act::D;FABPI:::bin::D;TRBM:::ind::D;BCL2:::mod::D|CP3A4:::sub::D;D6RB81:::sub::D;UD2B7:::sub::D;UD2B4:::sub::D;UD19:::sub::D;UD13:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D|S22A6:::inh:5.1:DC;S22AB:::inh::D;S22A8:::inh::D;SO1A2:::inh::D;MRP1:::inh::D;MRP4:::inh::D;MDR1:::sub::D;SO2B1:::sub::D|ALBU:::bin::D
Novobiocin|ok_inv_vet|GYRB::STAAU:inh:8.:DC;GYRB::STRPN::7.43:C;GYRB::MYCSM::7.34:C;GYRB::MYCS2::7.34:C;GYRB::ECOLI::7.1:C;TOP1::STAAU:inh::D||SO2B1:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;S22AB:::inh::D;S22A8:::inh::D;S22A6:::inh::D|
Benzylpenicillin|ok_vet|BLAT::ECOLX:::D;PBP3::STAA3:inh::D||SO1B1:::sub::D;SO3A1:::sub::D;SO4A1:::sub::D;SO2B1:::sub::D;S22AB:::inh::D;S22A4:::inh::D;S22A6:::inh::D;S22A5:::inh::D;S15A2:::inh::DC;S15A1:::inh::DC;S22A8:::inh::DC|
Nitrendipine|ok_inv|CAC1C:::inh:9.82:DC;CP2C9::::6.52:C;CP2CJ::::5.52:C;TRPA1::MOUSE::5.42:C;LMNA::::5.4:C;AA3R::::5.08:C;AA1R::RAT::5.05:C;GEMI::::5.:C;KCNH2::::5.:C;CAC1H:::inh::D;CA2D2:::inh::D;CAC1S:::inh::D;CAC1D:::inh::D;CCG1:::inh::D;CACB2:::inh::D;CA2D1:::inh::D|CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|ABCBB:::sub::D;MDR1:::inh::D|
Tocainide|ok|SCN5A:::inh::D|CP1A2:::inh::D||ALBU
Echothiophate|ok|CHLE:::inh::D|||ALBU
Praziquantel|ok_inv_vet|BLM::::8.49:C;P53::::6.9:C;NPSR1::::5.2:C;Schistosome_calcium_ion_Ca2_channels::Schistosoma:::D|CP3A7:::sub::D;CP3A5:::sub::D;CP343:::sub::D;CP2CJ:::sub::D;CP1A2:::sub::D;CP3A4:::sub::D||
Norfloxacin|ok|GBRP::RAT::7.7:C;GYRB::ECOLI::6.22:C;KDM4E::::5.9:C;CP2J2::::5.59:C;PGDH::::5.55:C;PARC::STAAU::5.46:C;HD::::5.45:C;NPSR1::::5.3:C;LMNA::::5.1:C;AL1A1::::5.05:C;TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A1:::inh::D;CP3A4:::inh::D;CP1A2:::inh::D|S22A6:::inh::D;S22A5:::inh::D|
Amoxicillin|ok_vet|PBPA::CLOPE:inh::D||S22A6:::inh::D;S15A2:::inh::D;S15A1:::inh::D|
Azlocillin|ok|PBPA::CLOPE:inh::D|||
Oxybutynin|ok_inv|ACM4::::9.56:C;ACM3:::ant:9.24:DC;ACM1:::ant:9.07:DC;ACM3::RAT::9.02:C;ACM5::::8.64:C;ACM1::RAT::8.23:C;ACM2::RAT::8.16:C;ACM2:::ant:8.09:DC;SGMR1::::7.99:C;SC6A3::::7.17:C;DRD3::::6.84:C;5HT2B::::6.3:C;CP2CJ::::6.22:C;SC6A2::::5.59:C|CP3A5:::sub::D;CP2D6:::inh::D;CP2C8:::inh::D;CP3A4:::inh::D||ALBU:::bin::D;A1AG1:::bin::D
Acetophenazine|ok|ANDR::RAT::6.1:C;ANDR;DRD1:::ant::D;DRD2:::ant::D|||
Isoprenaline|ok_inv|ADRB1:::ago:10.08:DC;ADRB2::CANLF::10.:C;ADRB2::RAT::10.:C;ADRB2:::ago:9.8:DC;ADRB3:::ago:9.01:DC;ADA1A::::8.82:C;ADRB1::RAT::8.28:C;ADRB3::RAT::7.89:C;ADRB2::CAVPO::7.75:C;ADRB2::BOVIN::6.96:C;ADRB1::MOUSE::6.66:C;LOX15::RABIT::5.75:C;DRD4::::5.54:C;DRD3::::5.33:C;TAU::::5.1:C;SODC;CAMP_phosphodiesterase::TRYCR:act::D;P55G:::ago::D;P85B:::ago::D;P85A:::ago::D;MK01:::ind::D|CP1A1:::inh::D||
Melatonin|ok_nutra_vet|MTR1A:::ago:10.77:DC;MTR1B:::ago:10.16:DC;MTR1C::XENLA::10.1:C;MTR1C::CHICK::9.75:C;MTR1B::CHICK::9.15:C;BLM::::8.8:C;NQO2::::7.56:DC;ACM1::RAT::7.2:C;CP2D6::::5.:C;CALR;PERE:::inh::D;CALM1;RORB:::ago::D;ESR1:::ant::D|CP1A2:::sub:5.3:DC;CP19A:::inh::D;I23O1:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP1B1:::inh::D;CP1A1:::inh::D;ASMT:::sub::DC;PERM:::inh::DC|S22A8:::inh::D|
Cefditoren|ok_inv|PBP2::STRR6:inh::D;PBPA::CLOPE:inh::D|||
Glipizide|ok_inv|NFKB1::::7.95:C;LMNA::::7.05:C;TSHR::::5.4:C;CP3A4::::5.13:C;PPARG:::ago::D;ABCC8:::inh::D|CP2C9:::sub:5.1:DC;UD11:::sub::D|ABCBB:::sub::D|ALBU:::bin::D
Clonazepam|ok_ill|GBRA2::BOVIN::9.07:C;GBRA1::::9.07:C;GBRP::RAT::8.77:C;NR1I2:::pag::D;TSPO;GABAR:::aga::D|ARY2:::sub::D;CP2E1:::inh::D;CP3A4:::sub::D||ALBU
Promethazine|ok_inv|HRH1:::ant:9.48:DC;ACM4:::ant:8.98:DC;ACM1:::ant:8.48:DC;ACM5:::ant:8.48:DC;ACM3:::ant:8.38:DC;5HT2C::::8.19:C;ACM2:::ant:7.92:DC;5HT2A:::ant:7.72:DC;ADA1B::RAT::7.68:C;ADA2B::::7.62:C;ADA1A::RAT::7.49:C;5HT2B::::7.37:C;LMNA::::7.25:C;ADA1D::::7.05:C;DRD2:::ant:7.:DC;SGMR1::::6.92:C;DRD3::::6.72:C;ADA2A::::6.59:C;ADA2C::::6.45:C;5HT6R::::5.95:C;HRH2:::ant:5.94:DC;DRD1::::5.86:C;5HT1A::RAT::5.83:C;SC6A4::::5.67:C;SC6A2::::5.38:C;SCN1A::::5.16:C;PRIO::::5.1:C;CALM1:::inh::D;ADA1A|CP2C9:::inh::D;CP2B6:::sub::D;CP2D6:::inh::D|MDR1:::inh::D|
Dihydrotachysterol|ok|VDR:::ago::D|||
Mequitazine|exp|HRH1:::ant::D|CP3A4:::inh::D;CP2D6:::sub::D||
Atazanavir|ok_inv|Pol_polyprotein::9HIV1:inh::D|CP1A2:::inh::D;CP2C8:::inh::D;UD11:::inh::D;CP2C9:::inh::D;CP3A4:::inh::D|SO1B3:::inh:6.43:DC;SO1B1:::inh:5.89:DC;SO2B1:::inh:5.29:DC;ABCBB:::sub::D;MRP1:::inh::D;MDR1:::inh::D|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Fludarabine|ok|AA1R::RAT::8.23:C;AA2AR::RAT::7.55:C;HIF1A::::5.2:C;DCK:::ago::D;DNA:::destbz::D;DPOLA:::inh::D;RIR1:::inh::D||S28A3;S29A1:::sub::D|
Perhexiline|ok_inv|ADA1B::RAT::6.7:C;ACM4::::6.3:C;ACM1::::6.19:C;ACM3::::6.18:C;ACM5::::6.1:C;SGMR1::::5.96:C;EGFR::::5.83:C;SC6A2::::5.49:C;FYN::::5.39:C;KCNH2::::5.11:DC;CPT2:::inh::D;CPT1A:::inh::D|CP2D6:::inh:6.03:DC;CP3A4:::sub::D;CP2B6:::sub::D||
Diphenhydramine|ok_inv|HRH1::CAVPO::9.:C;HRH1:::ant:7.83:DC;ACM4::::7.28:C;TPO::::7.2:C;ACM1::::7.08:C;ACM5::::6.94:C;ACM3::::6.86:C;ACM1::RAT::6.7:C;ACM2:::ant:6.43:DC;5HT2A::::6.43:C;5HT2C::::6.29:C;5HT2B::::6.15:C;KCNH2::::5.59:C;SC6A2::::5.45:C;SCN1A::::5.22:C|CP2D6:::inh:5.4:DC;PGH1:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D|S22A5:::inh::D;S22A2:::inh::D|
Atorvastatin|ok|HMDH:::inh:9.64:DC;HMDH::RAT::8.42:C;CYSP::TRYCR::5.15:C;NR1I3:::lig::D;HDAC2:::inh::D;AHR:::ago::D;DPP4:::inh::D|CP3A4:::sub:5.29:DC;UD13:::sub::D;UD11:::sub::D;CP2B6:::ind::D;CP2CJ:::inh::D;CP2C9:::inh::D;CP2D6:::inh::D;CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D|SO1B1:::inh:6.22:DC;ABCBB:::sub::D;MRP2:::sub::D;SO1B3:::sub::D;SO2B1:::sub::D;MRP1:::sub::D;MRP5:::sub::D;MRP4:::sub::D;SO1A2:::sub::D;MDR1:::inh::D|ALBU:::bin::D
Etidronic_acid|ok|LMNA::::5.9:C;VATA:::inh::D;PTPRS:::inh::D;Hydroxylapatite:::ant::D;Adenosine_triphosphate_ATP:::inh::D|||
Deslanoside|ok|TAU::::7.1:C;AT1A1:::inh::D|||
Tegaserod|ok_out|5HT4R:::ant_pago:9.:DC;5HT4R::CAVPO::8.2:C;5HT3A::::5.6:C;5HT2A:::ant::D;5HT2C:::ant::D;5HT2B:::ant::D|CP2E1:::inh::D;CP2D6:::inh::D;CP2C8:::inh::D;CP1A2:::inh::D|MDR1:::sub::D;ABCG2:::sub::D;SC6A4:::inh::D|
Vigabatrin|ok|GABT:::inh::D;GABR1:::ago::D|CP2C9:::ind::D|S36A1|
Diphenoxylate|ok_ill|KCNA3::::5.3:C;OPRD:::ago::D;OPRM:::ago::D|||
Streptomycin|ok_vet|PADI4;16S_ribosomal_RNA::Gut_flora:inh::D;RS12::ECOLI:inh::D||S22A6:::inh::D|
Orlistat|ok_inv|DGLA::::9.:C;FAAH1::RAT::8.:C;LIPP::PIG::7.92:C;ABHD6::::7.88:C;DGLA::MOUSE::7.7:C;ABHGA::::7.52:C;PAFA::::7.3:C;DGLB::::7.22:C;ABD12::::7.1:C;FAS:::inh:6.55:DC;NR1I2::::5.8:C;MEN1::::5.7:C;CNR1::::5.6:C;LIPG:::inh::D;LIPP:::inh::D|PA24A:::inh::D;CP3A4:::ind::D||
Emedastine|ok|HRH1::CAVPO::8.21:C;HRH1:::ant::D|||
Pilocarpine|ok_inv|ACM1:::ago:7.76:DC;ACM1::RAT::7.17:C;CP2AD::::5.85:C;ACM1::DROME::5.55:C;ACM1::MOUSE::5.16:C;ACM2::RAT::5.06:C;ACM4:::pag::D;ACM2:::ago::D;ACM3:::ago::D|CP2A6:::inh:5.52:DC;CP3A4:::inh::D||
Benzocaine|ok_inv|CP1A2::::5.7:C;RORG::MOUSE::5.15:C;LMNA::::5.1:C;SCNAA:::inh::D|EST1:::inh::D|MDR1:::inh::D|
Primaquine|ok|SC6A4::::8.08:C;NQO2:::inh:5.12:DC;K2C7;Fe_II_protoporphyrin_IX::PLAFA:ant::D|CP1A2:::sub_ind:6.74:DC;CP1B1:::ind::D;CP1A1:::ind::D;CP2D6:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Iloprost|ok_inv|PI2R:::ago:8.32:DC;PD2R2:::ago::D;TPA;PDE4D:::ind::D;PDE4C:::ind::D;PDE4B:::ind::D;PDE4A:::ind::D;PE2R1:::ago::D||SO3A1:::sub::D;SO2A1:::sub::D;SO2B1:::sub::D|
Deserpidine|ok|RORG::MOUSE::5.15:C;MEN1::::5.1:C;VMAT2:::inh::D|||
Pentolinium|ok|ACHB4:::ant::D;ACHA3:::ant::D;ACH10:::ant::D|||
Butenafine|ok|CP2D6::::6.52:C;SC6A4::::6.12:C;ADA2A::::5.86:C;SGMR1::::5.78:C;SC6A2::::5.41:C;ACES::::5.16:C;ERG1:::inh::D|||
Ouabain|ok|LMNA::::7.5:C;P53::::7.3:C;GEMI::::6.95:C;KLF5::::6.78:C;STAT3::::5.94:C;AT1A1:::inh:5.22:DC;AT1A3:::inh::D;AT1A2:::inh::D||SO1B1:::inh::D;SO1C1:::sub::D;SO1B3:::sub::D;SO4C1:::sub::D;S22A8:::inh::D;SO1A2:::inh::D|
Dimethyl_sulfoxide|ok_vet||CP3A4:::inh::D;CP2D6:::inh::D;CP2CJ:::inh::D||TTHY
Fluvastatin|ok|HDAC2:::inh::D;HMDH:::inh::D|CP2B6:::ind::D;UD2B7:::sub::D;UD13:::sub::D;UD11:::sub::D;CP2D6:::sub::D;CP2CJ:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;CP3A5:::sub::D;CP3A4:::inh::D;CP1A1:::sub_ind::D|MRP2:::sub::D;S15A1:::inh::D;SO2B1;SO1B3:::sub::D;SO1B1:::inh::D|
Oxamniquine|ok|DNA|CP2D6:::inh::D||
Leflunomide|ok_inv|LMNA::::8.49:C;PYRD::RAT::8.05:C;PYRD::MOUSE::7.52:C;NPSR1::::7.1:C;HD::::6.5:C;NPC1::::6.25:C;CP3A4::::6.2:C;RAB9A::::6.14:C;LUCI::PHOPY::6.05:C;SC6A3::::5.64:C;GEMI::::5.5:C;SC6A2::::5.34:C;SMN::::5.15:C;TPO::::5.1:C;ACM1::RAT::5.05:C;P53::::5.:C;PYRD:::inh:5.:DC;FAK2:::ant::D;AHR:::ago::D|CP1A2:::sub:7.2:DC;CP2C9:::inh::D|ABCG2:::sub::D|
Rosuvastatin|ok|HMDH:::inh:9.05:DC;HMDH::RAT::8.68:C;PDE6D::::5.9:C;ITAL:::inh_allo::D|CP2C9:::sub::D|NTCP;S22A8:::inh::D;MRP2:::sub::D;ABCG2:::sub::D;ABCBB:::sub::D;XCT;SO2B1;SO1B3;SO1B1:::inh::D;SO1A2;MRP4:::sub::D|ALBU:::sub::D
Flucytosine|ok_inv|TYSY::CANAL:inh::D;DNMT1;DNA:::cov::D|||
Pimozide|ok|DRD5::RAT::9.4:C;5HT7R::RAT::9.3:C;DRD2::BOVIN::9.22:C;KCNH2:::inh:8.52:DC;IMPA1::RAT::8.1:C;DRD2:::ant:7.93:DC;CAC1G::::7.4:C;SCN1A::::7.27:C;MK01::::7.2:C;5HT6R::::7.15:C;CAC1C::::6.79:C;SCN2A::RAT::6.47:C;OPRM::::6.43:C;OPRK::::6.:C;HIF1A::::5.9:C;GLRA1::::5.77:C;KCNK2::::5.74:C;UBP1::::5.7:C;MEN1::::5.55:C;FRIL::HORSE::5.5:C;OPRD::::5.42:C;MDR1A::MOUSE::5.31:C;LMNA::::5.25:C;NPSR1::::5.2:C;TAU::::5.2:C;ACM1::RAT::5.05:C;TPO::::5.:C;END4::ECOLI::5.:C;CP2CJ::::5.:C;CALM1:::inh::D;DRD3:::ant::D|CP3A4:::inh:5.5:DC;CP2D6:::inh:5.5:DC;CP1A2:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|MDR1:::inh:6.1:DC|
Capecitabine|ok_inv|RNA:::destbz::D;DNA:::destbz::D;TYSY:::inh::D|CP2C9:::inh::D;CDD:::sub::D;DPYD:::sub::D;EST1:::sub::D;TYPH:::sub::D||
Arbutamine|ok|ADRB1:::ago::D;ADRB2:::ago::D;ADRB3:::ago::D|||
Quinacrine|inv|ACM3::::6.58:C;RBP::CHICK::6.58:C;ACM4::::6.56:C;PRIO::::6.52:C;ACM2::::6.46:C;ACM1::::6.44:C;DRD3::::6.35:C;ADA2C::::6.25:C;5HT2A::::6.12:C;ADA2B::::6.08:C;ADA2A::::6.07:C;ADA1D::::5.99:C;ADA1B::RAT::5.72:C;ACM5::::5.57:C;ACES::::5.57:C;SC6A2::::5.54:C;SCN1A::::5.48:C;AOXA::::5.48:C;HRH2::::5.46:C;CHLE::HORSE::5.35:C;CAC1C::RAT::5.28:C;CAC1C::CAVPO::5.25:C;AOXA::RABIT::5.:C;PLCL1:::inh::D;PA24A:::inh::D;PLPL9:::inh::D;DNA:::itc::D|CP3A5:::sub::D;CP3A4:::sub::D;HNMT:::inh::D|MDR1:::inh::D;S22A2:::inh::D|
Sertraline|ok|SC6A4:::inh:10.12:DC;SC6A4::RAT::9.07:C;SC6A3:::inh:7.6:DC;SGMR1::::7.53:C;SC6A3::RAT::7.11:C;ADA2B::::7.08:C;ADA2A::::6.97:C;ACM1::::6.51:C;ADA1B::RAT::6.48:C;ACM4::::6.44:C;ACM5::::6.44:C;SC6A2:::idw:6.38:DC;5HT2C::::6.25:C;ADA2C::::6.19:C;5HT2A::::6.11:C;ACM2::::6.01:C;5HT2B::::5.67:C;CAC1C::RAT::5.64:C;MEN1::::5.45:C;MC5R::::5.37:C;KCNH2::::5.17:C;KMT2A::::5.1:C;S29A4;PGRC1,SGMR1:::inh:,7.53:DC|CP2CJ:::inh:6.51:DC;CP3A4:::sub:6.1:DC;CP2D6:::inh:5.85:DC;CP2E1:::sub::D;Q14097:::ind::D;AOFA:::sub::D;AOFB:::sub::D;CP2B6:::inh::D;CP2C9:::inh::D|MDR1:::inh::D|ALBU:::bin::D
Sibutramine|ok_ill_inv_out|SC6A3:::inh:6.3:DC;ADA2B::::5.96:C;SC6A4:::inh:5.96:DC;SC6A2:::inh:5.25:DC|CP3A4:::sub::D||
Levocabastine|ok_inv|NTR2::RAT::7.55:C;NTR2:::antp::D;HRH1:::ant::D|||
Methyprylon|ok_ill_out|GBRA1:::ago::D;GABAR:::aga::D|||
Trilostane|ok_inv_vet_out|ESR2:::alo::D;ESR1:::alo::D;3BHS2:::inh::D;3BHS1:::inh::D|CP3A4:::sub::D||
Heparin|ok_inv|ANT3:::pot::D;FA10:::inh::D;LYAM3:::inh::D;FGFR4;FGF4;FGF19;FGFR1;FGF1;FGFR2;FGF2;PLF4;HGF|HPSE:::sub::D||THBG:::sub::D
Miconazole|ok_inv_vet|LMNA::::8.05:C;CP121::MYCTU::7.14:C;CP51::MYCTU::6.7:C;CP17A::::6.61:C;THAS::::6.58:C;CP19A::RAT::6.4:C;SC6A4::::6.38:C;ACM4::::6.35:C;CP2J2::::6.24:C;ACM3::::6.18:C;ACM1::::6.02:C;DRD3::::5.96:C;5HT2A::::5.95:C;OPRD::::5.92:C;CP1A2::::5.9:C;SC6A3::::5.87:C;ADA2A::::5.83:C;ADA1D::::5.82:C;ACM2::::5.81:C;AA3R::::5.8:C;NK2R::::5.79:C;ADA2B::::5.78:C;MDR1B::MOUSE::5.7:C;OPRM::::5.61:C;OPRK::::5.58:C;5HT2C::::5.56:C;SC6A2::::5.54:C;CAC1C::RAT::5.52:C;DRD1::::5.51:C;5HT2B::::5.45:C;NK1R::::5.43:C;I23O1::::5.42:C;ADRB3::::5.39:C;FYN::::5.38:C;DRD2::::5.38:C;ANDR::RAT::5.33:C;5HT6R::::5.3:C;DRD4::::5.27:C;GRM6::::5.19:C;HRH2::::5.18:C;5HT1A::RAT::5.18:C;I23O2::MOUSE::5.17:C;AA1R::::5.14:C;ADRB1::::5.14:C;AGTR2::::5.11:C;MDR1A::MOUSE::5.11:C;AA2AR::::5.1:C;5HT1B::RAT::5.03:C;NR1I2:::pag::D;KCNH7:::inh::D;KCNH6:::inh::D;KCNH2:::inh::D;KCNN3:::inh::D;KCNN2:::inh::D;KCNN1:::inh::D;KCNN4:::inh::D;KCMB4:::inh::D;KCMB3:::inh::D;KCMB2:::inh::D;KCMB1:::inh::D;KCMA1:::inh::D;NOS2:::inh::D;NOS3:::inh::D;CP51::CANAL:inh::D|CP2CJ:::inh:7.8:DC;CP3A4:::inh:7.:DC;CP2C9:::inh:6.7:DC;CP51A:::inh:6.7:DC;CP19A:::inh:6.22:DC;CP2D6:::inh:6.:DC;C11B1:::inh::D;CP2E1:::inh::D;CP2B6:::inh::D;CP2A6:::inh::D|MDR1:::inh:5.7:DC|
Colistimethate|ok_vet|Bacterial_outer_membrane::Bacteria:destbz::D|||
Cefuroxime|ok|PBPA::CLOPE:inh::D||S15A2:::inh::D;S15A1:::inh::D|
Papaverine|ok_inv|RORG::MOUSE::8.55:C;PDE10:::inh:7.77:DC;PDE10::RAT::7.44:C;ACM1::RAT::7.25:C;PDE3A::::6.55:C;PDE3B::::6.38:C;CBP::::6.25:C;CP2CJ::::6.12:C;ADRB1::RAT::6.:C;LMNA::::5.7:C;CP3A4::::5.7:C;PDE2A::::5.64:C;HIF1A::::5.6:C;FFP::BACIU::5.55:C;TSHR::::5.5:C;PDE4A::::5.18:C;LOX12::::5.15:C;KCNH2::::5.14:C;MK01::::5.1:C;PDE5A::::5.06:C;PDE1B::BOVIN::5.06:C;PDE1A::::5.05:C;NFKB1::::5.:C;CP2D6::::5.:C;ADA1B::RAT::5.:C;CP1A2::::5.:C;PDE4B:::inh::D|||
Chlorpheniramine|ok|HRH1:::ant:9.04:DC;HRH1::RAT::8.7:C;HRH1::CAVPO::8.06:C;KCNH2::::5.96:C;SCN1A::::5.:C;SC6A3:::inh::D;SC6A2:::inh::D;SC6A4:::inh::D|CP3A5:::sub::D;CP2D6:::inh::D;CP3A4:::sub::D;CP3A7:::sub::D|S22A1:::inh::D;S22A2:::inh::D|
Nifedipine|ok|CAC1C:::inh:9.4:DC;CAC1C::RABIT::9.:C;CAC1D::RAT::8.92:C;CAC1C::RAT::8.85:C;CAC1C::CAVPO::8.59:C;TSHR::::6.8:C;AMPC::ECOLI::6.45:C;TRPA1::MOUSE::6.4:C;HIF1A::::6.3:C;CCR2::::6.07:C;CAC1B::::5.95:C;LMNA::::5.95:C;CHLE::HORSE::5.92:C;CAC1D:::inh:5.87:DC;I23O2::MOUSE::5.82:C;TPO::::5.8:C;MYLK::::5.69:C;AA1R::RAT::5.54:C;CP2J2::::5.51:C;RORG::MOUSE::5.5:C;TAU::::5.45:C;BLM::::5.4:C;ACES::ELEEL::5.4:C;AA3R::::5.39:C;CP2C9::::5.39:C;AA1R::::5.35:C;CP2CJ::::5.27:C;SMN::::5.25:C;KCNA5::::5.21:C;PLIN5::::5.15:C;AL1A1::::5.1:C;HCD2::::5.1:C;5HT2C::::5.02:C;ABHD5::::5.02:C;NR1I2;CAC1H:::inh::D;KCNA1:::inh::D;CALM1:::inh::D;CAC1S:::inh::D;CA2D1:::inh::D;CACB2:::inh::D|CP1A2:::inh:7.4:DC;CP3A4:::duo:5.25:DC;CP2B6:::ind::D;CP1A1:::inh::D;CP2E1:::inh::D;CP2D6:::inh::D;CP2C8:::inh::D;CP2A6:::sub::D|ABCBB:::sub::D;SO1B1:::inh::D;MRP2:::ind::D;MDR1:::duo::D;MRP3:::ind::D|
Trimethaphan|ok_inv|ACHA::TETCF::5.15:C;ACH10:::ant::D|CHLE:::sub::D||
Atovaquone|ok|PYRD::RAT::6.15:C;PYRD:::inh::D;PYRD::PLAF7:inh::D;CYB::PLAFA:inh::D|CP3A4:::sub::D;CP2C9:::inh::D|MDR1:::inh::D|
Amiodarone|ok_inv|SGMR1::::9.:C;EBP::::7.6:C;KCNH2:::inh:7.52:DC;ERG2::YEAST::7.21:C;ADA2A::::6.93:C;5HT2C::::6.67:C;CAC1C::::6.57:C;DRD3::::6.39:C;ACM4::::6.3:C;5HT2B::::6.23:C;THB::::6.22:DC;ACM1::::6.2:C;THA::::6.19:DC;ACM3::::6.17:C;FFP::BACIU::6.15:C;FYN::::6.09:C;5HT2A::::5.99:C;ACM5::::5.97:C;SC6A4::::5.91:C;SO1A4::RAT::5.74:C;ACM2::::5.74:C;SC6A3::::5.7:C;MDR1A::MOUSE::5.68:C;SC6A2::::5.65:C;OPRD::::5.55:C;LEF::BACAN::5.46:C;NFKB1::::5.45:C;CCR2::::5.37:C;DRD1::::5.34:C;SCN1A::::5.32:C;AL1A1::::5.3:C;ADA2B::::5.23:C;DRD4::::5.21:C;TSHR::::5.2:C;NK2R::::5.19:C;DRD2::::5.18:C;OPRK::::5.18:C;OPRM::::5.11:C;BKRB2::::5.11:C;FDFT::::5.1:C;MC5R::::5.05:C;5HT6R::::5.04:C;ERBB2::::5.04:C;P53::::5.:C;AA3R::::5.:C;MK01::::5.:C;PPARG:::ago::D;CA2D2:::inh::D;CAC1H:::inh::D;ADRB1:::ant::D|CP2C9:::inh:8.1:DC;CP2C8:::sub:5.82:DC;CP1A2:::inh:5.5:DC;CP3A4:::inh:5.2:DC;CP2J2:::inh::D;CP2A6:::inh::D;CP1A1:::sub::D;CP2CJ:::inh::D;CP2D6:::inh::D|MDR1:::duo:5.49:DC;S22A2:::inh::D;ABCBB:::inh::D|
Diazoxide|ok|LMNA::::6.95:C;CP1A2::::5.7:C;THB::::5.2:C;CP2D6::::5.1:C;KCJ11:::ind:5.06:DC;S12A3;KCMA1;AT1A1;CAH2:::inh::D;CAH1:::inh::D|GLNA:::inh::D||
Gliclazide|ok|VEGFA;ABCC8:::bin::D|CP2CJ:::sub::D;CP2C9:::sub::D||ALBU
Phenacemide|ok|SCN1A:::inh::D|||
Ambenonium|ok|ACES::BOVIN::9.92:C;ACES:::inh::D|CHLE:::inh::D||
Proflavine|ok|MEN1::::6.45:C;TetR_family_transcriptional_regulator::MYCSM:::D;QACR::STAAU:::D;THRB;DNA:::itc::D|||
Tolbutamide|ok_inv|ACM1::RAT::7.55:C;LMNA::::6.65:C;LEF::BACAN::5.4:C;ALBU::RAT::5.1:C;KCNJ1:::inh::D;ABCC8:::inh::D|CP2CI:::sub::D;CP2CJ:::sub::D;CP2C8:::inh::D;CP2C9:::sub::D|SO2B1:::sub::D;S15A2:::inh::D;S22A6:::inh::D;SO1A2:::inh::D;S15A1:::inh::D|ALBU::::5.22:DC
Anisindione|ok|SMN::::5.4:C;RAB9A::::5.35:C;PGDH::::5.35:C;NPC1::::5.25:C;LOX5::RAT::5.04:C;P53::::5.:C;VKGC:::inh::D|||
Dutasteride|ok_inv|GLRA1::::6.48:C;S5A1:::inh::D;S5A2:::inh::D|CP3A5:::sub::D|VMAT2::MOUSE:bin::D;SC6A3::MOUSE:bin::D|A1AG1:::bin::D;ALBU:::bin::D
Econazole|ok|THAS::::7.54:C;CP2CJ::::7.4:C;CP51A::::7.3:C;CP121::MYCTU::7.14:C;CP2C9::::6.7:C;CP51::MYCTU::6.7:C;SC6A4::::6.65:C;ACM4::::6.53:C;CP1A2::::6.52:C;CP17A::::6.49:C;ACM3::::6.42:C;CP2D6::::6.4:C;OPRD::::6.29:C;ACM1::::6.2:C;SC6A3::::6.18:C;ACM2::::5.94:C;5HT2A::::5.94:C;HRH2::::5.81:C;ADA2A::::5.79:C;DRD3::::5.79:C;AA3R::::5.74:C;NK2R::::5.7:C;OPRM::::5.64:C;SC6A2::::5.62:C;ADA2B::::5.57:C;DRD4::::5.49:C;OPRK::::5.46:C;DRD2::::5.37:C;ADA1D::::5.36:C;5HT2B::::5.36:C;ADRB3::::5.34:C;DRD1::::5.34:C;5HT6R::::5.3:C;5HT2C::::5.2:C;NK1R::::5.19:C;ANDR::RAT::5.17:C;MMP9::::5.16:C;ADRB1::::5.13:C;I23O2::MOUSE::5.12:C;AA2AR::::5.09:C;I23O1::::5.09:C;ADA1A::RAT::5.07:C;SGMR1::::5.05:C;5HT1A::RAT::5.03:C;AA1R::::5.01:C;5HT1B::RAT::5.:C;NR1I2:::pag::D;CP51::CANAL:ant::D|CP3A4:::inh:7.3:DC;CP2E1:::inh::D;CP19A:::inh::D||
Bicalutamide|ok|ANDR::RAT::7.85:C;ANDR:::ant:7.72:DC;ANDR::MOUSE::6.17:C;PRGR::::5.74:C;PRGR::RABIT::5.25:C;PRGR::RAT::5.14:C|CP2D6:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D;CP3A4:::inh::D||
Rabeprazole|ok_inv|LMNA::::7.55:C;DRD3::::6.1:C;ADA2B::::6.1:C;AA3R::::5.74:C;FAS::::5.23:C;AL1A1::::5.22:C;TAU::::5.:C;ATP4A:::inh::D|CP2C8:::inh::D;CP2D6:::inh::D;CP2C9:::inh::D;CP1A2:::ind::D;CP1A1:::ind::D;CP2CJ:::inh::D;CP3A4:::inh::D|ABCG2:::inh::D|
Prednicarbate|ok_inv|GCR:::ago::D|CP3A4:::sub_ind::D||
Proguanil|ok|LMNA::::5.7:C;CP1A2::::5.1:C;DRTS::PLAFK:inh::D;DYR:::inh::D|CP2D6:::inh:5.:DC;CP2C9:::sub::D;CP2CJ:::sub::D||
Pioglitazone|ok_inv|PPARG:::ago:7.06:DC;CAH2::::6.94:C;AOFB::::6.7:DC;ABCBB::::6.52:C;CISD1::::6.43:C;PPARG::MOUSE::6.26:C;PPARG::RAT::6.15:C;CISD1::RAT::6.:C;ABCBB::RAT::5.7:C;AOFB::RAT::5.68:C;PPARA::::5.18:DC;PPARD|CP2C9:::sub::D;PGH1:::sub::D;CP3A4:::sub_ind::D;CP2C8:::inh::D|SO1B1:::inh::D;SO1B3:::inh::D|
Tiludronic_acid|ok_inv_vet|MMP2::::5.14:C;PTN1:::inh::D;VATA:::inh::D;Hydroxylapatite:::ant::D;Adenosine_triphosphate_ATP:::inh::D|||
Doxacurium|ok|ACHA2:::ant::D;ACM2:::ant::D|CHLE:::sub::D||
Carvedilol|ok_inv|ADRB1:::ant:9.99:DC;ADRB2:::ant:9.78:DC;ADRB1::RAT::9.09:C;ADA1D:::ant:9.05:DC;ADA1B::RAT::8.71:C;ADRB3::::8.51:C;ADA1A::RAT::8.5:C;5HT1A::RAT::8.5:C;ADA2C:::ant:7.89:DC;5HT2B::::7.82:C;ADA2A:::ant:7.4:DC;ADA2B:::ant:7.37:DC;DRD2::::7.31:C;5HT2C::::7.22:C;5HT2A::::6.93:C;SC6A4::::6.93:C;5HT4R::CAVPO::6.74:C;DRD3::::6.71:C;KCNH2:::inh:6.46:DC;SC6A2::::6.27:C;5HT1B::RAT::6.23:C;SC6A3::::6.17:C;5HT6R::::6.15:C;DRD1::::6.13:C;RORG::MOUSE::6.:C;KCNK2::::5.8:C;CAC1C::RABIT::5.44:C;S22A2::::5.12:C;KCNKA::::5.12:C;KCNJ2:::inh::D;KCNJ4:::inh::D;HIF1A:::mod::D;LYAM2:::inh::D;ADA1B:::ant::D;VCAM1:::inh::D;CXA1;ANFB;VEGFA;NDUC2:::inh::D;ADA1A:::ant::D|UD2B7:::sub::D;UD2B4:::sub::D;UD11:::sub::D;CP2E1:::sub::D;CP1A1:::sub::D;CP3A4:::sub::D;CP1A2:::sub::D;CP2D6:::sub::D;CP2C9:::sub::D;XDH:::inh::D|MDR1:::inh:5.34:DC|ALBU:::bin::D
Levofloxacin|ok_inv|STRP::STRP1::5.81:C;TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP2C9:::inh::D;CP3A4:::inh::D;CP1A2:::inh::D|S47A2:::inh::D;S47A1:::inh::D;S22A4:::inh::D;S22A2:::inh::D;S22A6:::sub::D;MDR1:::inh::D|
Sulfinpyrazone|ok|AL1A1::::6.1:C;MEN1::::5.6:C;HCD2::::5.3:C;FPR1::::5.:C;PGDH::::5.:C;KDM4E::::5.:C;NR1I2:::act::D;S22AC:::inh::D|CP3A4:::sub_ind:5.2:DC;CP2C9:::inh:5.:DC;CP2C8:::inh::D;CP2B6:::ind::D|ABCBB:::sub::D;MRP6:::inh::D;MRP5:::inh::D;MRP4:::inh::D;MRP3:::inh::D;MRP1:::inh::DC;MRP2:::inh::DC|FABPI
Cefapirin|ok_vet|PBPA::CLOPE:inh::D|||
Cefadroxil|ok_vet_out|S15A2::RAT::5.52:C;PBP2::STRR6:inh::D;PBP1B::STRR6:inh::D;PBPA::STRR6:inh::D;PBP3::STREE:inh::D||S15A2:::inh:5.6:DC;S22A6:::inh:5.21:DC;S22A8:::inh:5.06:DC;S22A5:::inh::D;S15A1:::inh::D|
Micafungin|ok_inv|FKS1::ASPNC:inh::D|ARSA:::sub::D;COMT:::sub::D||
Doxepin|ok_inv|HRH1:::ant:9.6:DC;KCNH2:::inh:5.19:DC;HRH4:::bin::D;5HT6R:::bin::D;5HT1A:::ant::D;ADA1D:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;5HT2C:::ant::D;5HT2B:::ant::D;5HT2A:::ant::D;SC6A4:::inh::D;SC6A2:::inh::D;HRH2:::ant::D|CP3A4:::sub::D;CP1A2:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP2D6:::inh::D|MDR1:::sub::D|A1AG1:::bin::D;ALBU:::bin::D
Amifostine|ok_inv|ACM1::RAT::7.95:C;DRD3::::6.18:C;ENPP1:::ind::D;PPBN:::ind::D|PPBT:::sub::D||
Diclofenamide|ok_inv|CAH7:::inh:8.22:DC;CAH2:::inh:8.1:DC;CAH5B::::7.68:C;CAH13::::7.64:C;CAH13::MOUSE::7.64:C;CAH1:::inh:7.6:DC;CAH9::::7.47:C;CAN::CANAL::7.42:C;CAH12::::7.3:C;CAH6::::7.1:C;CAH5A::::7.09:C;CAH15::MOUSE::7.02:C;CAH4:::inh:7.02:DC;CAN::YEAST::6.99:C;CAH::METTE::6.82:C;CAH14::::6.46:C;LMNA::::6.45:C;CYNT::HELPY::6.44:C;CAH4::BOVIN::6.42:C;MTCA1::MYCTU::6.06:C;MTCA2::MYCTU::5.7:C;CAH3:::inh::D|||
Sulfoxone|ok|Dihydropteroate_synthetase::PLAFA:inh::D|||
Diphenylpyraline|ok_inv|SC6A3::RAT::6.38:C;CP2D6::::5.2:C;SC6A3:::inh::D;HRH1:::ant::D|||
Cloxacillin|ok_inv_vet|DACA::ECOL6:inh::D;Cell_division_protein::PSEAI:inh::D;PBP2::STRPN:inh::D;PBP2A::STRR6:inh::D;AMPC::ECOLI:ind::D;PBPA::CLOPE:inh::D||S22A6:::inh::D;S15A2:::inh::D;S15A1:::inh::D|ALBU
Flavoxate|ok|LMNA::::5.9:C;CP1A2::::5.2:C;CP2D6::::5.1:C;CP3A4::::5.:C;ACM1:::ant::D;ACM2:::ant::D|||
Nefazodone|ok_out|5HT2A:::ant:8.24:DC;SC6A4::RAT::6.86:C;5HT1A:::ant:6.8:DC;SC6A4:::inh:6.7:DC;SC6A2:::inh:6.44:DC;SC6A3:::inh:6.44:DC;SC6A3::RAT::5.62:C;MEN1::::5.5:C;KCNH2:::ant::D;ADA1A:::ant::D;ADA2A:::ant::D;ADA1B;5HT2C:::ant::D|CP3A4,CP343,CP3A5,CP3A7:::inh:7.82,,,:DC;CP3A4:::inh:7.82:DC;CP2D6:::inh::D;Q14097:::inh::D|ABCBB:::sub:5.38:DC;MDR1:::duo:5.33:DC;SO2B1:::inh::D;SO1B3:::inh::D|
Cefprozil|ok|PBPA::STRPN:inh::D;PBPX::STRPN:inh::D;PBP2::STRPN:inh::D|||
Desipramine|ok_inv|ADA1A::RAT::9.6:C;SC6A3::::9.31:C;SC6A2:::inh:9.22:DC;HRH1::RAT::9.1:C;SC6A4:::inh:7.7:DC;5HT2A:::ant:6.8:DC;SC6A4::RAT::6.79:C;ACM1::RAT::6.5:C;5HT3A::RAT::6.46:C;KCNH2::::5.86:C;SCN5A::::5.82:C;SC6A2::MOUSE::5.8:C;CAC1C::CAVPO::5.77:C;SCN1A::::5.62:C;S22A1::RAT::5.55:C;HRH2::CAVPO::5.42:C;SC6A3::RAT::5.19:C;SC6A4::MOUSE::5.03:C;NFKB1::::5.:C;S22A2::RAT::5.:C;ADA2A,ADA2B,ADA2C:::bin::D;DRD2:::bin::D;5HT2C:::bin::D;5HT1A:::bin::D;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;ADA1A,ADA1B,ADA1D:::ant::D;HRH1:::ant::D;ASM:::inh::D;ADRB1;ADRB2:::ant::D|CP2D6:::inh:5.4:DC;CP2E1:::inh::D;CP2B6:::inh::D;CP3A4:::inh::D;CP1A2:::sub::D|S22A1:::inh:5.27:DC;S22A4:::inh::D;S22A5:::inh::D;S22A2:::inh::D;S22A3:::inh::D;MDR1:::inh::D|A1AG1
Candicidin|ok_out|Ergosterol::CANAL:ant::D|CP3A4:::inh::D||
Sertaconazole|ok_inv|I23O1::::5.08:C;CP51::CANAL:inh::D|||
Thiamylal|ok_vet|GBRA1:::ago::D;KCNJ8:::inh::D;KCJ11:::inh::D|CP2C9:::sub::D;CP3A4:::sub_ind::D;CP2E1:::sub::D||
Gemifloxacin|ok_inv|PARC::STAAU::6.52:C;GYRB::ECOLI::6.3:C;GYRB::STAAU::5.25:C;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A2:::inh::D||
Bupropion|ok|ACHA::::8.1:C;ACHB2::::7.92:C;ACHB4::::7.82:C;SC6A3::RAT::6.43:C;SC6A3:::inh:6.36:DC;SC6A2:::inh:6.35:DC;CP2CJ::::5.7:C;ACHA7::::5.1:C;5HT3A:::neg::D;ACHA3:::ant::D|CP2E1:::sub::D;CP2C9:::sub::D;CP2D6:::inh::D;CP2B6:::sub::D|S22A2:::inh::D|A1AG1:::ant::D
Trimetrexate|ok_inv|DYR::MOUSE::10.22:C;DYR::PNECA::9.15:C;DYR:::inh:8.85:DC;DYR::CANAX::8.72:C;DYR::RAT::8.52:C;DRTS::TOXGO::8.29:C;DRTS::TRYCR::8.18:C;DYR::ECOLI::8.:C;DYR::LACCA::7.57:C;DYR::YEAST::7.38:C|||
Bretylium|ok|AT1A1:::inh::D|||
Halothane|ok_vet|GABAR:::aga::D;NPSR1;GBG2;GBRA1;AT2C1;ATPD;KCNN4:::inh::D;NU1M:::inh::D;KCNJ3:::inh::D;KCNJ6:::inh::D;OPSD;GLRA1:::alo::D;NMDE1:::ant::D;NMD3B:::ant::D;NMD3A:::ant::D;KCMA1:::inh::D;KCNK9:::bin::D;KCNK3:::bin::D|CP2C9:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;CP3A4:::sub::D;CP2E1:::sub::D||ALBU
Dinoprost_tromethamine|ok_vet|LMNA::::8.:C;PI2R:::ant::D;PF2R:::ago::D||SO3A1;SO2A1;S22AB;S22A8;S22A7;S22A6;S22A2|
Chloroprocaine|ok|SCNAA:::inh::D;NMD3A:::ant::D;ACH10:::ant::D;5HT3A:::ant::D;SC6A3:::inh::D|CHLE:::sub::D||
Terazosin|ok|ADA1B::RAT::10.99:C;ADA1A:::ant:10.4:DC;ADA1A::RAT::10.15:C;ADA1A::BOVIN::9.9:C;ADA1D::RAT::9.77:C;ADA1D:::ant:9.7:DC;OPRM::RAT::9.7:C;ADA1B:::ant:9.68:DC;5HT1D::::9.48:C;CASB::RAT::9.44:C;ADA2C::RAT::9.4:C;ADA1B::MESAU::9.16:C;AA3R::::9.07:C;ADA1A::RABIT::8.3:C;ADA2B::RAT::8.11:C;NQO2::::8.11:C;ADA2B::::7.89:C;ADA2B::MOUSE::7.89:C;ADA2C::::7.62:C;ADA2A::::7.47:C;ADA2A::BOVIN::6.97:C;LMNA::::6.95:C;KDM4E::::6.2:C;5HT2A::RAT::5.82:C;KCNH2:::inh:5.8:DC;S47A1::::5.8:C;ADA2A::RAT::5.78:C;S22A1::::5.74:C;5HT1A::RAT::5.63:C;5HT2B::::5.58:C;SMN::::5.4:C;MMP1::::5.39:C;ADA2A::PIG::5.39:C;HD::::5.35:C;CP3A4::::5.2:C;MMP9::::5.16:C;LEF::BACAN::5.1:C;DRD4::::5.08:C;SCN1A::::5.:C;TGFB1:::ind::D;KCNH7:::inh::D;KCNH6:::inh::D||MDR1:::inh::D|
Amdinocillin|inv_out|PBP1B::STRR6:inh::D;PBP2::STRR6:inh::D;PBPA::STRR6:inh::D;PBP3::STREE:inh::D;MRDA::ECOLI:inh::D;PBP2A::STRR6:inh::D|||
Calcium_chloride|ok|S10AD|||
Ofloxacin|ok|STE24::YEAST::5.71:C;PGDH::::5.5:C;KDM4E::::5.5:C;STRP::STRP1::5.43:C;TRYP::PIG::5.03:C;HCD2::::5.:C;TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A2:::inh::D|ABCBB:::sub::D;S22A4:::inh::D;MRP2:::inh::D;S22A6:::inh::D;MRP1:::inh::D;S22A5:::inh::D|
Cilostazol|ok_inv|BLM::::7.:C;PDE3A:::inh:6.72:DC;RORG::MOUSE::5.5:C;MK01::::5.45:C;AL1A1::::5.1:C;CP2C9::::5.:C|CP3A4:::sub:5.:DC;CP2D6:::sub::D;CP1A2:::sub::D;CP2CJ:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D||
Itraconazole|ok_inv|CXCR1::::7.:C;MDR1A::MOUSE::6.7:C;CCR4::::6.7:C;MDR1B::MOUSE::6.15:C;V2R::::6.1:C;CYSP::TRYCR::5.52:C;CP51A:::inh:5.44:DC;FYN::::5.41:C;CP51::CANGA:inh::D|CP3A4:::inh:7.15:DC;CP2E1:::inh::D;CP1A1:::ind::D;CP2B6:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D|MDR1:::inh:7.52:DC;SO2B1:::inh::D|
Procarbazine|ok_inv|CP1A2::::5.8:C;LMNA::::5.5:C;CP2CJ::::5.3:C;LOX15::::5.1:C;AOFA,AOFB:::inh::D;DNA:::cov::D|XDH:::sub::D||
Arsenic_trioxide|ok_inv|LMNA::::5.15:C;PML;HDAC1;CDN1A;AKT1:::ind::D;MK01:::ind::D;MK03:::ind::D;CCND1:::ant::D;JUN:::ind::D;TRXR1:::inh::D;IKKB:::ind::D|CP3A4:::inh::D|MDR1:::sub::D;MRP2:::ind::D|ALBU:::sub::D
Guanethidine|ok|LMNA::::5.85:C;SC6A2:::ind::D|||
Moclobemide|ok_inv|AOFA,AOFB:::ant:8.3,5.97:DC;AOFA::RAT::8.3:C;AOFB::RAT::5.97:C;5HT1A::::5.3:C|AOFA:::inh:8.3:DC;AOFB:::inh:5.97:DC;CP2C9:::sub::D;CP2D6:::inh::D;CP2CJ:::inh::D||
Kanamycin|ok_inv_vet|FABH::ECOLI::5.17:C;16S_ribosomal_RNA::Gut_flora:inh::D;RS12::ECOLI:inh::D|KKA1::ECOLX:sub::D;KANU::STAAU:sub::D;AAC2::MYCTU:sub::D||
Orphenadrine|ok|ACM4::::7.77:C;ACM5::::7.7:C;ACM1::::7.44:C;ACM3::::7.43:C;5HT2A::::6.9:C;ACM2::::6.87:C;HRH1:::ant:6.84:DC;HRH1::RAT::6.79:C;SC6A4::::6.61:C;5HT2C::::6.55:C;5HT6R::::6.28:C;ADA2A::::6.09:C;KCNH2::::6.07:C;ADA2B::::6.06:C;5HT2B::::5.67:C;S22A2::::5.6:C;SC6A2:::inh:5.58:DC;NMDZ1:::ant:5.22:DC;HRH2::::5.16:C;SCNAA:::inh::D;NMD3A:::ant::D;NMD3B:::ant::D;NMDE4:::ant::D|CP2D6:::inh:6.4:DC;CP1A2:::inh::D;CP2E1:::inh::D;CP3A4:::inh::D;CP2B6:::inh::D||
Phenobarbital|ok_inv|SCN2A::RAT::5.6:C;NR1I2:::act::D;NMDA:::ant::D;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA1:::pot::D|UD2B7:::ind::D;UD11:::ind::D;CP4B1:::ind::D;CP3A7:::ind::D;CP2CI:::sub::D;CP1A1:::ind::D;CP3A5:::ind::D;CP2E1:::sub_ind::D;CP2A6:::ind::D;CP1A2:::ind::D;CP3A4:::ind::D;CP2C8:::ind::D;CP2B6:::ind::D;CP2C9:::sub_ind::D;CP2CJ:::sub_ind::D|MRP2:::ind::D;SO2A1:::ind::D;MRP1:::ind::D;ABCBB:::ind::D;MRP3:::ind::D;MDR1:::sub_ind::D|
Escitalopram|ok|SC6A4::RAT::9.05:C;SC6A4:::inh:9.:DC;NFKB1::::5.95:C;CP2C9::::5.5:C;LOX15::::5.2:C;ACM1::RAT::5.2:C;SC6A3::RAT::5.09:C;SC6A3:::inh::D;SC6A2:::inh::D;DRD2:::inh::D;ADA2A,ADA2B,ADA2C:::inh::D;5HT2C:::inh::D;ADA1A,ADA1B,ADA1D:::inh::D;5HT2A:::inh::D;5HT1A:::inh::D;HRH1:::inh::D;ACM1:::inh::D|CP3A4:::sub:6.:DC;CP2CJ:::sub:5.5:DC;AOFA,AOFB:::sub::D;CP2D6:::inh::D|MDR1:::sub::D|
Cyclizine|ok|HRH1:::ant:8.35:DC;5HT2A::::7.19:C;ACM4::::6.92:C;ACM3::::6.8:C;ACM1::::6.79:C;5HT2B::::6.62:C;ACM2::::6.39:C;ACM5::::6.34:C;5HT2C::::6.27:C;ADA2A::::6.24:C;ADA1D::::6.22:C;SC6A3::::6.22:C;DRD3::::5.99:C;ADA1B::RAT::5.86:C;CP2D6::::5.21:C;RORG::MOUSE::5.2:C;ST1E1:::inh::D|CP2C9:::inh::D||
Idarubicin|ok|LMNA::::6.6:C;MTOR::::6.38:C;PMP22::::6.37:C;HD::::6.2:C;MEN1::::5.75:C;TAU::::5.45:C;TOP2A:::inh::D;DNA:::itc::D|CP2D6:::sub::D;CP2C9:::sub::D|MRP1:::inh::D|
Chlormezanone|ok_out|LMNA::::5.25:C;TSPO:::ago::D|||
Podofilox|ok|GCR::::7.85:C;HIF1A::::7.8:C;LMNA::::7.55:C;TBB::PIG::6.46:C;TBB4B::::6.46:C;TBB2B::BOVIN::6.34:C;TBA1A::PIG::6.34:C;CP3A4::::6.22:C;LEF::BACAN::6.1:C;VE2::HPV1::5.98:C;NR0B1::::5.67:C;CP2C9::::5.4:C;CP2CJ::::5.3:C;TBB5:::inh::D;TBA4A:::inh::D;TOP2A:::inh::D|||
Rescinnamine|ok|ACE:::inh::D|||
Ifosfamide|ok|LMNA::::7.25:C;MEN1::::5.55:C;NR1I2;DNA|PGH1:::sub::D;CP2CI:::sub::D;CP2A6:::sub::D;CP2C8:::sub_ind::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP3A5:::sub::D;CP3A4:::duo::D;CP2B6:::sub::D||
Propafenone|ok|ADRB2:::ant:7.44:DC;5HT2B::::7.24:C;5HT2A::::6.73:C;5HT2C::::6.7:C;ADRB1:::ant:6.69:DC;ADRB3::::6.5:C;KCNH2:::inh:6.36:DC;5HT6R::::6.06:C;5HT1A::RAT::6.03:C;SGMR1::::5.96:C;SCN5A:::inh:5.92:DC;ADA1B::RAT::5.85:C;SC6A3::::5.83:C;CAC1C::CAVPO::5.74:C;KCJ11::::5.66:C;ADA1A::RAT::5.6:C;SC6A2::::5.52:C;KCNK3::::5.29:C;KCNK2::::5.12:C|CP1A2:::inh:5.48:DC;CP2D6:::inh:5.34:DC;CP3A4:::sub::D|MDR1:::inh:6.49:DC|
Naloxone|ok_vet|OPRM:::ant:9.66:DC;OPRK:::ant:9.6:DC;OPRM::RAT::9.4:C;OPRM::CAVPO::9.17:C;OPRK::RAT::9.:C;SGMR1::RAT::9.:C;AA3R::::8.8:C;OPRD::RAT::8.6:C;OPRK::CAVPO::8.51:C;OPRM::BOVIN::8.3:C;OPRM::MOUSE::7.99:C;CCR5::MOUSE::7.98:C;OPRD:::ant:7.72:DC;OPRD::MOUSE::7.35:C;OPRK::MOUSE::6.9:C;CP2D6::::5.7:C;EST1;TLR4:::inh::D;ESR1:::ant::D;CREB1|UD11:::sub::D;CP3A4:::inh::D|MDR1:::sub::D;SO1A2:::inh::D|ALBU:::sub::D
Domperidone|ok_inv_vet|DRD2::RAT::9.28:C;DRD2:::ant:9.05:DC;DRD3::RAT::8.99:C;DRD3:::ant:8.46:DC;5HT2A::::7.96:C;KCNH2::::7.24:C;ADA1B::RAT::7.06:C;ADA1A::RAT::6.94:C;NFKB1::::6.85:C;ADA2C::::6.83:C;HRH1::::6.81:C;ADA1D::::6.28:C;5HT2C::::6.16:C;ADA2B::::6.01:C;ADA2A::::5.99:C;AOXA::::5.92:C;SC6A4::::5.79:C;5HT2B::::5.78:C;OPRM::::5.77:C;S47A1::::5.64:C;HIF1A::::5.6:C;SC6A2::::5.59:C;OPRK::::5.55:C;LMNA::::5.25:C;S22A2::::5.1:C|CP2D6:::sub:5.5:DC;CP1A2:::sub:5.2:DC;CP2C8:::sub::D;CP2B6:::sub::D;CP3A4:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|MDR1:::sub::D|
Fluoxymesterone|ok_ill|ANDR:::ago:9.52:DC;DHI2:::inh::D;GCR:::ant::D;PRLR:::ant::D;ESR1:::ant::D|||SHBG:::ant::D
Pergolide|ok_inv_vet_out|DRD2:::ago:9.45:DC;DRD3:::ago:9.07:DC;DRD2::RAT::9.:C;DRD5::RAT::8.8:C;5HT1A:::ago:8.74:DC;DRD3::RAT::8.62:C;5HT2A:::ago:8.41:DC;DRD2:S194A:RAT::8.4:C;5HT1A::RAT::8.07:C;DRD1::BOVIN::7.74:C;5HT6R::::7.74:C;ADA2B:::ago:7.54:DC;DRD2:S197A:RAT::7.4:C;5HT1B::RAT::7.4:C;ADA2C::RAT::7.39:C;ADA2A::BOVIN::7.39:C;DRD2::BOVIN::7.32:C;5HT2B:::ago:7.31:DC;ADA2A:::ago:7.:DC;KCNH2::::6.92:C;5HT3A::RAT::6.85:C;5HT2C:::ago:6.7:DC;ADA2C:::ago:6.69:DC;DRD1:::ago:6.47:DC;ADA1B::RAT::6.26:C;ADA1D:::ago:6.13:DC;ADA1A::RAT::6.11:C;ADA1B:::ago::D;ADA1A:::ago::D;5HT1B:::ago::D;DRD5:::ago::D;5HT1D:::ago::D;DRD4:::ago::D|CP2D6:::inh:6.7:DC;CP3A4:::inh::D||
Iophendylate|ok||||
Ciclopirox|ok_inv|AT1A1:::bin::D|||
Desflurane|ok|GABAR:::aga::D;GLRA1:::ago::D;GRIA1:::ant::D;KCNA1:::ind::D;AT2C1:::inh::D;ATPD;NU1M|||ALBU
Clindamycin|ok_vet|23S_ribosomal_RNA::Gut_flora:inh::D;RL10::SHIFL:inh::D|CP3A4:::inh::D||
Dexfenfluramine|ok_ill_inv_out|SGMR1::::6.66:C;5HT1A::RAT::5.71:C;5HT2C:::ago::D;SC6A4:::inh::D|CP2E1:::inh::D;CP1A2:::sub::D;CP2D6:::inh::D||
Oxymorphone|ok_inv_vet|SGMR1::RAT::10.89:C;OPRM::CAVPO::9.27:C;OPRM::RAT::9.01:C;OPRM::MOUSE::8.33:C;OPRD:::ant:7.35:DC;OPRK::CAVPO::7.24:C;OPRD::RAT::7.09:C;OPRK::::7.05:C;OPRK::RAT::7.02:C;OPRD::MOUSE::6.21:C;OPRM:::ago::D|CP2D6:::sub::D;CP3A4:::sub::D||
Acebutolol|ok_inv|ADRB1:::pag:6.37:DC;5HT1A::RAT::5.:C;ADRB2:::pag::D|CP2D6:::inh::D|MDR1:::sub::D|
Brinzolamide|ok|CAH2:::inh:10.05:DC;CAH6::::9.05:C;CAH7::::8.55:C;CAH12::::8.52:C;CAH1:::inh:8.52:DC;CAN::CANAL::8.52:C;CAH13::MOUSE::8.:C;CAH13::::7.96:C;CAH14::::7.62:C;CAH5B::::7.52:C;CAH9::::7.44:C;CAH4::BOVIN::7.35:C;CAH4:::inh:7.34:DC;CAH5A:::inh:7.3:DC;CAH15::MOUSE::7.21:C;CAN::YEAST::6.94:C;MTCA2::MYCTU::6.9:C;CYNT::HELPY::6.68:C;MTCA1::MYCTU::6.08:C;CAH3:::inh::D|CP3A4:::sub::D||
Flecainide|ok_out|LMNA::::5.9:C;KCNH2:::inh:5.41:DC;SCN5A:::inh:5.19:DC;KCND2::RAT::5.:C;RYR2:::inh::D;SCN4A:::inh::D|CP2C9:::inh::D;CP1A2:::sub::D;CP2D6:::inh::D|S47A1:::inh::D;MDR1:::sub::D|ALBU:::bin::D;A1AG1,A1AG2:::bin::D
Estramustine|ok_inv|RECQ1::::5.09:C;ESR2;ESR1:::ago::D;MAP1A:::ant::D;MTAP2:::ant::D|CP3A4:::sub::D|MDR1:::inh::D|
Captopril|ok|ACE:::inh:9.92:DC;ACE::RABIT::8.77:C;RENI::::8.77:C;ACE::RAT::8.7:C;THRB::::7.32:C;LKHA4:::inh:7.15:DC;DAPE::HAEIN::5.74:C;BKRB1;MMP9:::inh::D;MMP2:::inh::D||S22A6:::inh::D;S15A1:::inh::D;MDR1:::inh::D|ALBU
Zopiclone|ok|GBRP::RAT::7.54:C;TAU::::6.05:C;RECQ1::::5.85:C;TSPO:::ago::D;GBRA5:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2E1:::sub::D;PGH1:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP3A4:::sub::D||
Tubocurarine|ok|S47A1::::5.03:C;ACHA7;ACES:::inh::D;5HT3A:::ant::D;ACHA2:::ant::D|CHLE:::sub::D|S22A2;S22A1:::sub::D|
Bromocriptine|ok_inv|DRD3:::ago:9.69:DC;DRD2:::ago:9.3:DC;5HT2A:::ago:8.75:DC;ADA1B::RAT::8.71:C;ADA1A::RAT::8.55:C;5HT1A::RAT::8.49:C;DRD2:S197A:RAT::8.4:C;5HT2B:::ago:8.28:DC;ADA2A:::ago:8.26:DC;DRD2::RAT::8.1:C;DRD2:S194A:RAT::8.1:C;5HT6R::::8.:C;ADA1D:::ago:7.82:DC;ADA2B:::ago:7.8:DC;5HT1A:::ago:7.62:DC;DRD5::RAT::7.55:C;5HT1B::RAT::7.33:C;ADA2C:::ago:7.12:DC;5HT2C:::ago:6.56:DC;ADA2C::RAT::6.29:C;ADA2A::BOVIN::6.29:C;ADRB1::::5.86:C;DRD1:::ago:5.84:DC;ANDR::RAT::5.82:C;RORG::MOUSE::5.45:C;TAU::::5.4:C;LMNA::::5.3:C;MDR1B::MOUSE::5.19:C;MDR1A::MOUSE::5.13:C;5HT7R:::ant::D;ADA1B:::duo::D;ADA1A:::duo::D;DRD5:::ago::D;5HT1B:::ago::D;DRD4:::ant::D;5HT1D:::ago::D|CP3A4:::inh:5.7:DC|MDR1:::inh:5.55:DC|
Rifapentine|ok_inv|RPOC::MYCTU:inh::D|CP3A4,CP343,CP3A5,CP3A7:::ind::D;CP2B6:::ind::D;CP2CJ:::ind::D;CP2C8:::ind::D;CP3A4:::sub_ind::D;CP2C9:::ind::D||
Levetiracetam|ok|CAC1B:::inh::D;SV2A:::ago::D||MDR1:::sub::D|
Nadolol|ok|RECQ1::::6.9:C;ADRB2:::ant::D;ADRB1:::ant::D||S47A2:::sub::D;S47A1:::sub::D;PO2F2:::sub::D;PO2F1:::sub::D;MDR1:::sub::D|A1AG1,A1AG2:::bin::D
Mitoxantrone|ok_inv|TPO::::7.6:C;LMNA::::7.15:C;ACM2::::7.11:C;ACM4::::7.05:C;MTOR::::6.83:C;ACM1::::6.74:C;S47A1::::6.72:C;S47A2::::6.28:C;CSK2B::::6.18:C;BTK::::6.:C;FYN::::5.9:C;DYR1A::RAT::5.9:C;LOX15::RABIT::5.75:C;5HT2C::::5.73:C;NFKB1::::5.7:C;P53::::5.7:C;ERBB2::::5.69:C;NSD2::::5.63:C;KCNH2::::5.53:C;SO1B3::::5.51:C;MK01::::5.4:C;SC6A2::::5.31:C;ACM1::RAT::5.3:C;TOP2A:::inh:5.28:DC;EGFR::::5.27:C;HIF1A::::5.1:C;IMPA1::RAT::5.:C;HD::::5.:C;DNA:::itc::D|CP3A4:::inh::D;CP1B1:::inh::D;CP2E1:::sub_ind::D|MRP1:::inh:8.82:DC;ABCG2:::sub::D;MDR1:::duo::D|
Flumazenil|ok|GBRA2::BOVIN::10.05:C;GBRG2:::ant:9.35:DC;GBRG2::RAT::9.3:C;GBRA5:::ant:9.3:DC;GBRP::RAT::9.1:C;GBRA1:::ant:9.1:DC;GBRA4::::8.7:C;GBRB2::::8.24:C;TSHR::::7.5:C;RORG::MOUSE::7.:C;CP2CJ::::5.8:C;ACM1::RAT::5.55:C;END4::ECOLI::5.:C;GABAR:::aga::D|||
Lomustine|ok_inv|STMN4:::ant::D;DNA:::cov::D|CP2D6:::inh::D;CP3A4:::inh::D||
Sparfloxacin|ok_out|MK01::::5.35:C;TOP2A:::inh::D;GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D|CP1A2:::inh::D|MDR1:::sub::D;MRP2:::inh::D;S22A5:::inh::D|
Dezocine|ok_inv|OPRM:::ago:7.42:DC;OPRK:::ant::D|||
Levobunolol|ok|ADRB2:::ant:9.26:DC;ADRB1:::ant:8.4:DC;ADRB3::::6.59:C;SGMR1::::6.49:C;5HT1A::RAT::5.78:C;SC6A4::::5.58:C;TSHR::::5.1:C|CP2D6:::sub::D||
Clarithromycin|ok|SO1B1::::5.51:DC;SO1B3::::5.48:DC;MK01::::5.4:C;KCNH2;RL10::SHIFL:inh::D|CP3A4:::inh:5.26:DC;CP3A5:::inh::D|MDR1:::inh:5.42:DC;ABCBB:::sub::D;S22A7:::inh::D|
Ceftriaxone|ok|OXDA::::5.:C;PBP2::STRR6:inh::D|GLNA:::ind::D|S22A6:::inh:6.64:DC;S22AB:::inh:5.62:DC;S22A8:::inh:5.36:DC;S15A2:::inh::D;S15A1:::inh::DC|ALBU
Fomepizole|ok_vet|ADH1E::HORSE::7.89:C;CATA:::inh::D;ADH1G:::inh::D;ADH1B:::inh::D;ADH1A:::inh::D|CP2A6:::inh::D;CP2E1:::sub_ind::D||
Metipranolol|ok|ADRB1:::ant::D;ADRB2:::ant::D|CP2D6:::sub::D||
Estazolam|ok_ill|GABAR:::aga::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRA5:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP3A4:::sub::D||
Finasteride|ok|S5A2:::inh:9.74:DC;S5A2::RAT::9.55:C;BLM::::8.55:C;S5A1::RAT::8.38:C;S5A1:::inh:7.58:DC;CP2CJ::::6.:C;CP2C9::::5.7:C;RORG::MOUSE::5.4:C;LMNA::::5.25:C;MK01::::5.2:C;TPO::::5.:C;AK1D1:::inh::D|CP3A4:::sub:5.7:DC;CP3A7:::sub::D;CP3A5:::sub::D|S12A5::MOUSE:mod::D|
Anastrozole|ok_inv|CP19A:::inh:9.89:DC|UD14:::sub:5.33:DC;CP2C9:::inh::D;CP1A2:::inh::D;UD2B7:::sub::D;UD13:::sub::D;CP2C8:::inh::D;CP3A5:::sub::D;CP3A4:::inh::D|MDR1:::sub::D|
Halofantrine|ok|KCNH2:::inh:7.4:DC;CAC1C::::5.72:C;PLM2::PLAFA:inh::D;Fe_II_protoporphyrin_IX::PLAFA:ant::D|CP2C8:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D;CP2D6:::inh::D||
Dantrolene|ok_inv|CISD1::::5.69:C;LMNA::::5.2:C;TAU::::5.:C;RYR1:::ant::D|||THBG:::sub::D
Rifaximin|ok_inv|NR1I2:::ago:5.66:DC;FRIL::HORSE::5.:C;RPOB::ECOLI:inh::D|CP2C8:::ind::D;CP2CJ:::ind::D;CP3A4:::sub_ind::D||
Ketamine|ok_vet|NMDZ1::::6.38:C;NMDZ1::RAT::6.21:C;CAC1C::::5.74:C;ACHA::TETCF::5.31:C;NOS1:::inh::D;CHLE:::inh::D;Alpha_7_nicotinic_cholinergic_receptor_subunit:::ant::D;5HT3A:::pot::D;5HT1A,5HT1B,5HT1D,5HT1E,5HT1F:::ant::D;5HT2A,5HT2B,5HT2C:::ant::D;ACM1,ACM2,ACM3,ACM4,ACM5:::bin::D;OPRM:::bin::D;OPRK:::ago::D;SC6A2:::inh::D;OPRD:::bin::D;DRD2:::ago::D;NK1R:::ant::D;NMD3A:::ant::D|CP2C8:::sub::D;PGH1:::sub::D;CP2B6:::sub::D;CP3A4:::sub_ind::D;CP2C9:::sub::D||
Budesonide|ok|GCR:::ant:8.69:DC;GCR::RAT::8.54:C;TPO::::8.:C;NFKB1::::7.25:C;ANDR::RAT::5.96:C;MMP9::::5.7:C;ANXA1:::sub::D|CP3A4,CP343,CP3A5,CP3A7:::sub_ind:5.1,,,:DC;CP3A4:::sub_ind:5.1:DC;CP2CJ:::ind::D;CP2C9:::ind::D;CP2C8:::ind::D;CP2B6:::ind::D;CP1B1:::ind::D;CP2A6:::ind::D;CP3A5:::ind::D|S22A8:::sub::D;SO1A2:::sub::D;MDR1:::sub::D;ABCBB:::sub::D|ALBU:::bin::D;CBG:::bin::D
Aminophylline|ok|LMNA::::6.:C;TAU::::5.1:C;HDAC2:::act::D;AA3R:::ant::D;AA1R:::ant::D;PDE3A:::inh::D|CP3A4:::sub::D;CP2E1:::sub::D;CP1A2:::sub::D||
Quetiapine|ok|ADA1A,ADA1B,ADA1D:::ant:8.35,7.,7.32:DC;ADA1A::::8.35:C;HRH1:::ant:8.34:DC;H10::::8.:C;ADA1B::RAT::7.9:C;5HT2A:::ant:7.47:DC;ADA1A::RAT::7.46:C;HRH1::RAT::7.4:C;HRH1::CAVPO::7.4:C;ADA2B:::ant:7.34:DC;ADA1D::::7.32:C;ACM1:::ant:7.25:DC;ADA2C:::ant:7.21:DC;5HT7R:::lig:7.2:DC;DRD2:::ant:7.2:DC;5HT1A:::ant_pago:7.1:DC;ADA2A:::ant:7.06:DC;ADA1B::::7.:C;ACM4:::lig:6.9:DC;5HT2B::::6.87:C;DRD2::RAT::6.74:C;DRD1:::ant:6.67:DC;5HT2A::RAT::6.66:C;5HT1A::RAT::6.64:C;DRD3:::lig:6.6:DC;SGMR1::::6.02:C;ACM3:::ant:5.99:DC;ACM2:::lig:5.92:DC;AMPC::ECOLI::5.85:C;5HT2C:::lig:5.85:DC;5HT6R:::ant:5.85:DC;DRD4:::lig:5.8:DC;ACM5:::lig:5.67:DC;KCNH2::::5.24:C;DRD5:::lig::D;5HT3A:::lig::D;5HT1E:::lig::D;5HT1D:::lig::D;5HT1B:::lig::D|CP3A7;CP2D6:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D;CP3A5:::sub::D|MDR1:::sub::D|
Enoxaparin|ok|ANT3:::pot::D;FA10:::inh::D|PERM:::inh::D||
Mivacurium|ok|CHLE;ACM3:::ant::D;ACM2:::ant_pago::D;ACHA2:::ant::D|||
Levacetylmethadol|ok_inv|KCNH2::::5.66:C;ACHA3:::ant::D;ACHB4;OPRM:::ago::D|CP3A4:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D||
Encainide|ok_out|SCN5A:::inh::D|CP2D6:::sub::D||
Paclitaxel|ok_vet|LMNA::::8.74:C;TBB3::::8.11:C;GEMI::::7.65:C;TBB4B::::7.51:C;ITB3::::7.47:C;PMP22::::7.32:C;MTOR::::6.88:C;SO1B1::::6.55:C;TBB::PIG::6.28:C;THB::::6.15:C;TBB2B::BOVIN::6.08:C;RORG::MOUSE::5.95:C;OPRD::::5.83:C;NK2R::::5.69:C;CCKAR::::5.64:C;MEN1::::5.35:C;MERTK::::5.31:C;CYSP::TRYCR::5.3:C;BXA1::CLOBO::5.28:C;FFP::BACIU::5.:C;NR1I2:::ind::D;TAU;MTAP2;MAP4;BCL2:::inh::D;TBB1:::inh::D|CP3A4:::sub_ind:5.9:DC;CP1B1:::inh::D;CP19A:::inh::D;CP2C8:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D|SO1B3:::sub:6.59:DC;MDR1:::inh:5.59:DC;MRP2:::sub::D;MRP7:::inh::D;MRP1:::inh::D;ABCBB:::inh::D|
Pemoline|ok_ill_inv_out|SC6A3::::6.38:C;RAB9A::::5.9:C|||
Diphenidol|ok_out|ACM4::::7.42:C;ACM3:::ant:7.28:DC;ACM1:::ant:7.11:DC;SGMR1::::6.97:C;CP2D6::::6.9:C;ACM2:::ant:6.56:DC;5HT2A::::6.13:C;DRD3::::6.11:C;ACM5::::6.07:C;DRD2::::5.96:C;ADA1B::RAT::5.58:C;SCN1A::::5.47:C|||
Saquinavir|ok_inv|CAC1C::::5.72:C;NK2R::::5.68:C;THAS::::5.66:C;5HT1A::RAT::5.61:C;OPRK::::5.56:C;OPRM::::5.41:C;DRD3::::5.28:C;V1AR::::5.15:C;S22A1::RAT::5.08:C;OPRD::::5.:C;Pol_polyprotein::9HIV1:inh::D|CP3A4:::inh:6.77:DC;CP2D6:::inh::D;CP2C8:::inh::D;CP3A5:::inh::D;CP3A7:::inh::D|MDR1:::duo:5.8:DC;ABCBB:::sub::D;SO2B1:::inh::D;MRP2:::sub::D;MRP1:::sub::D;SO1B1:::inh::D;ABCG2:::inh::D;SO1A2:::inh::D;S22A1:::inh::D|ALBU;A1AG1
Metoclopramide|ok_inv|5HT4R::CAVPO::8.24:C;LMNA::::8.15:C;DRD3::::7.8:C;ACM1::RAT::7.45:C;DRD2:::ant:7.38:DC;5HT3A:::ago:7.3:DC;DRD3::RAT::7.21:C;DRD2::BOVIN::7.1:C;DRD2::RAT::6.98:C;5HT3A::RAT::6.8:C;5HT3B::MOUSE::6.7:C;5HT2B::::6.4:C;5HT4R:::ago:6.1:DC;5HT4R::RAT::6.1:C;ADA2A::::5.99:C;5HT2A::::5.98:C;5HT2C::::5.9:C;5HT1B::RAT::5.11:C;ADA2C::RAT::5.11:C;ACM1:::ago::D|CP2D6:::inh:6.1:DC;CP1A2:::sub::D;CP3A4:::sub::D|MDR1:::sub::D|A1AG1:::bin::D
Dexamethasone|ok_inv_vet|GCR:::ago:9.7:DC;MCR::::9.44:C;TSHR::::7.9:C;GCR::RAT::7.66:C;PRGR::::6.36:C;ANDR::::5.85:C;NR1I2::RAT::5.59:C;NR1I2:::ago::D;NOS2:::neg::D;ANXA1:::ago::D;NR0B1:::sti::D|C11B1:::inh::D;CP4AB:::ind::D;CP343:::ind::D;CP2E1:::ind::D;CP2C8:::ind::D;CP2CJ:::ind::D;CP2B6:::ind::D;CP2A6:::ind::D;CP1A1:::duo::D;CP17A:::inh::D;CP3A7:::sub_ind::D;CP3A5:::sub_ind::D;DHI1:::sub::D;CP3A4:::duo::D;DHI2:::sub::D|SO1A2:::inh::D;ABCG2:::inh::D;MRP2:::ind::D;ABCBB:::ind::D;S22A8:::sub::D;MDR1:::duo::D|ALBU:::bin::D
Levodopa|ok|ACM1::RAT::7.15:C;HCD2::::6.5:C;TYDP1::::6.3:C;FYN::::5.67:C;LOX15::RABIT::5.65:C;EGFR::::5.54:C;LCK::::5.43:C;HIF1A::::5.:C;DRD4:::ago::D;DRD3:::ago::D;DRD2:::ago::D;DRD5:::ago::D;DRD1:::ago::D|DDC:::sub::D|LAT2;LAT1;MOT10:::inh::D;S15A1:::inh::D|ALBU:::bin::D
Sevoflurane|ok_vet|GABAR:::aga::D;NU1M;ATPD;AT2C1:::inh::D;KCNA1:::ind::D;GRIA1:::ant::D;GLRA1:::ago::D;GBRA1:::ago::D|CP3A4:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;CP2E1:::sub::D||ALBU
Bromodiphenhydramine|ok|HRH1:::ant::D||S22A6|
Aripiprazole|ok_inv|DRD2:::ant_pago:9.7:DC;5HT2B:::ANT:9.44:DC;5HT1A::RAT::9.4:C;5HT2A:::ant_pago:9.1:DC;DRD1::RAT::9.1:C;DRD2::RAT::9.1:C;DRD3:::ant_pago:9.:DC;5HT1A:::pag:8.25:DC;5HT2A::RAT::8.15:C;5HT7R:::ant_pago:7.99:DC;5HT2C:::ant_pago:7.66:DC;HRH1:::ant:7.6:DC;ADA1A:::ant:7.59:DC;5HT2C::RAT::7.59:C;H10::::7.55:C;SC6A4:::mod:7.5:DC;DRD3::RAT::7.42:C;DRD4:::ant_pago:7.24:DC;5HT6R:::ant:7.05:DC;HRH1::CAVPO::7.:C;5HT1D:::ant:7.:DC;ADA1B::RAT::7.:C;ADA1B:::ant:7.:DC;ADA2A:::ant:7.:DC;ADA2C:::ant:7.:DC;DRD1:::ant_pago:6.51:DC;5HT3A:::ant:6.3:DC;DRD4::RAT::6.29:C;KCNH2::::6.22:C;RORG::MOUSE::6.15:C;MDR1::::6.11:C;5HT5A:::lig:6.:DC;ADA2B:::ant:6.:DC;5HT1B:::ant:6.:DC;DRD5:::ant_pago:5.98:DC;SC6A4::RAT::5.97:C;LYAG::::5.75:C;SC6A3:::mod::D;NMDA:::lig::D;OPRD:::lig::D;OPRM:::lig::D;OPRK:::lig::D;ACM5:::lig::D;ACM4:::lig::D;ACM3:::lig::D;ACM2:::lig::D;ACM1:::lig::D;HRH4:::lig::D;HRH3:::lig::D;HRH2:::lig::D;ADRB2:::lig::D;ADRB1:::lig::D;5HT1E:::ant::D|CP2D6:::sub::D;CP3A5:::sub::D;CP3A7:::sub::D;CP3A4:::sub::D||ALBU:::bin::D
Chlorprothixene|ok_exp_inv_out|CP1A2::::5.8:C;CP2D6::::5.6:C;LEF::BACAN::5.4:C;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;HRH1:::ant::D;5HT2C:::ant::D;5HT2B:::ant::D;5HT2A:::ant::D;DRD3:::ant::D;DRD1:::ant::D;DRD2:::ant::D||MDR1:::inh::D|
Epoprostenol|ok|PTGIS:::ind::D;PI2R:::ago::D;P2Y12:::ago::D|||
Gemfibrozil|ok|TTHY::::7.:C;FABPL::RAT::5.73:C;SO1B1:::inh:5.39:DC;SMN::::5.35:C;SO1B3:::inh:5.15:DC;CISD1::::5.14:C;SO2B1:::inh::D;S22A8:::inh::D;PPARA:::ago::D|CP2C8:::inh:5.39:DC;CP2C9:::inh:5.2:DC;UDB17:::sub::D;UD2B4:::sub::D;UD19:::sub::D;UD13:::inh::D;UD11:::inh::D;UD2B7:::sub::D;CP3A4:::sub::D;CP1A2:::inh::D;CP2CJ:::inh::D||ALBU:::bin::D
Clomipramine|ok_inv_vet|ADA1A::RAT::10.4:C;SC6A4:::inh:10.33:DC;HRH1::RAT::9.7:C;5HT3A::RAT::8.3:C;5HT2B::RAT::8.08:C;HRH1::::8.01:C;ACM4::::7.89:C;5HT2C:::ant:7.74:DC;5HT2A:::ant:7.72:DC;SC6A4::RAT::7.7:C;ACM1::::7.66:C;ACM3::::7.44:C;ACM5::::7.42:C;ADA2B::::7.34:C;DRD3::::7.33:C;ADA2C::RAT::7.29:C;DRD2::RAT::7.25:C;SC6A2:::inh:7.19:DC;SC6A4::MOUSE::7.15:C;ADA1B::RAT::7.14:C;ACM2::::7.07:C;ADA1D::::7.06:C;ACM1::RAT::7.:C;5HT6R::::6.95:C;DRD2::::6.86:C;5HT2B:::ant:6.82:DC;ADA2C::::6.69:C;IMPA1::RAT::6.35:C;ADA2A::::6.28:C;DRD1::::6.25:C;SGMR1::::6.24:C;TSHR::::6.2:C;HRH2::CAVPO::6.14:C;SC6A2::MOUSE::6.05:C;SC6A3::RAT::6.:C;HRH2::::5.7:C;SC6A3::::5.66:C;TYTR::TRYBB::5.47:C;5HT1B::RAT::5.3:C;TYTR::TRYCR::5.19:C;GSTP1:::inh::D|CP2D6:::inh:5.7:DC;CP1A2:::sub:5.3:DC;CP3A4:::sub::D;CP2CJ:::sub::D|MDR1:::inh::D|ALBU:::sub::D
Chloroxine|ok|MKNK2::::7.92:C;RORG::MOUSE::7.1:C;STRP::STRP1::6.83:C;HCD2::::6.3:C;LOX12::::6.:C;HS90A::::5.98:C;LOX15::::5.8:C;HD::::5.55:C;P53::::5.5:C;LOX5::::5.44:C;LMNA::::5.4:C;OPRK::::5.34:C;AL1A1::::5.3:C|||
Bepridil|ok_out|KCNH2:::inh:7.64:DC;CAC1C::CAVPO::6.68:C;SCN1A::::6.08:C;CAC1C::::6.:C;SCN5A::::5.43:C;CP2C9::::5.37:C;LEF::BACAN::5.32:C;PDE1A:::inh::D;PDE1B:::inh::D;CALM1:::bin::D;TNNC1;KCNQ1:::inh::D;AT1A1:::inh::D;CA2D2:::inh::D;CAC1H:::inh::D;CAC1A:::inh::D|CP3A4:::sub::D;CP2D6:::inh::D|MDR1:::inh::D|
Decamethonium|ok|NFKB1::::6.2:C;HRH3::::6.09:C;ACES::MOUSE::5.46:C;ACES:::inh:5.23:DC;LMNA::::5.1:C;ACM1::RAT::5.05:C;ACHB2;ACHA4;ACHA2:::pag::D|CHLE:::inh::D||
Alimemazine|ok_vet|HRH1:::ant::D|||
Isocarboxazid|ok|LMNA::::5.5:C;AOFB:::inh::D;AOFA:::inh::D|||
Docetaxel|ok_inv|NR1I2:::bin::D;TAU;MAP4;MTAP2;BCL2;TBB1|CP1B1:::bin::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::inh::D|MRP1:::sub::D;MRP2:::sub::D;ABCG2:::sub::D;S22A7:::sub::D;SO1B3:::sub::D;MRP7:::sub::D;MDR1:::sub::D|
Iodixanol|ok||||
Olsalazine|ok|IFNG;TPMT:::inh::D|||
Gliquidone|ok_inv|LMNA::::5.85:C;HIF1A::::5.6:C;KDM4E::::5.1:C;CP3A4::::5.:C;KCNJ8:::inh::D;ABCC8:::inh::D|CP2C9:::sub::D||
Mitiglinide|inv|PPARG:::ago::D;ABCC8:::inh::D|UD2B7:::sub::D;UD13:::sub::D||
Ergometrine|ok|5HT2A::::9.2:C;5HT1B::RAT::8.89:C;5HT6R::::8.82:C;5HT2B::::8.58:C;5HT1A::RAT::8.33:C;5HT2C::::7.96:C;ADA2B::::6.88:C;DRD2::::6.74:C;DRD3::::6.71:C;ADA2A::::6.2:C;DRD1::::5.53:C;ADA1A:::ago::D|CP3A4:::sub::D|MDR1:::inh::D|
Dasatinib|ok_inv|ABL1:M351T:::10.8:DC;ABL1:F317L:::10.72:DC;ABL1:H396P:::10.6:DC;ABL1::::10.54:DC;ABL1:Q252H:::10.43:DC;EPHB6::::10.41:C;ABL1:F317I:::10.39:DC;ABL1:E255K:::10.33:DC;ABL1:Y253F:::10.24:DC;LCK::MOUSE::10.19:C;EPHA3::::10.03:C;ABL2::::9.77:DC;FYN::::9.7:DC;LCK::::9.7:DC;BLK::::9.68:C;SRC::::9.68:DC;EPHA5::::9.62:DC;EPHA8::::9.62:C;ABL1:G250E:::9.6:DC;YES:::inh:9.52:DC;TXK::::9.52:C;FRK::::9.51:DC;HCK::::9.5:C;EPHB4::::9.47:DC;EPHB2::::9.41:C;DDR2::::9.4:C;SRC::CHICK::9.4:C;EPHB1::::9.35:C;PGFRA::::9.33:C;DDR1::::9.3:C;FGR::::9.3:DC;KIT:L576P::ant:9.24:DC;LYN::::9.24:DC;CSF1R::::9.24:C;KIT:::ant:9.21:DC;SRMS::::9.2:C;PGFRB:::ant:9.2:DC;KIT:A829P::ant:9.18:DC;KIT:V559D::ant:9.17:DC;SIK2::::9.1:C;EPHA2:::ant:9.07:DC;CSK::::9.:DC;EPHA4::::8.92:C;BTK::::8.89:DC;BMX::::8.85:C;KIT:D816H::ant:8.8:DC;ACK1::::8.6:C;KIT:D816V::ant:8.59:DC;GAK::::8.59:C;KIT:V559D-V654A::ant:8.57:DC;MP2K5::::8.48:C;SIK1::::8.41:C;EPHA1::::8.39:C;PTK6::::8.3:C;EPHB3::::8.16:C;BLK::MOUSE::8.1:C;TNI3K::::7.96:C;TEC::::7.89:C;M4K5::::7.8:C;ERBB3::::7.74:C;EGFR::::7.7:C;MK14::::7.57:DC;SIK3::::7.55:C;RIPK2::::7.51:C;TESK1::::7.48:C;ERBB4::::7.4:C;M3K20::::7.35:DC;BMR1B::::7.28:C;TBA1A::RAT::7.26:C;MYT1::::7.2:C;ACVR1::::7.1:C;EGFR:G719S:::7.1:C;M3K19::::7.1:C;LIMK2::::7.07:C;MK13::::7.:C;TYK2::::6.96:C;EGFR:L861Q:::6.96:C;LIMK1::::6.94:C;ABL1:T315I:::6.92:DC;EGFR:L858R:::6.92:C;PMYT1::::6.89:C;M3K2::::6.85:C;ERBB2::::6.8:C;RAF1::::6.79:C;EGFR:G719C:::6.77:C;COQ8A::::6.72:C;KSYK::::6.7:C;WEE2::::6.7:C;AVR2A::::6.68:C;STK36::::6.68:C;TGFR1::::6.64:C;NLK::::6.59:C;M3K3::::6.55:C;M3K4::::6.51:C;ACV1B::::6.48:C;RET:M918T:::6.41:C;MK11::::6.39:C;MINK1::::6.37:C;RET::::6.36:C;ACVL1::::6.34:C;NEK11::::6.33:C;BRAF::::6.3:C;BRAF:V600E:::6.24:C;AVR2B::::6.24:C;MP2K1::::6.2:C;SLK::::6.2:C;JAK3::::6.19:C;M4K3::::6.19:C;CDPK1::PLAF7::6.19:C;STK35::::6.11:C;FGFR1::::6.06:C;M4K1::::6.01:C;TAOK1::::6.:C;JAK2::::6.:C;SBK1::::5.92:C;STK10::::5.92:C;MRCKG::::5.92:C;DYRK3::::5.9:C;AURKB::::5.9:C;VGFR2::::5.9:C;FGFR3::::5.9:C;DMPK::::5.89:C;M4K2::::5.89:C;MP2K2::::5.85:C;FGFR2::::5.85:C;KC1E::::5.82:C;E2AK4::::5.8:C;STK26::::5.72:C;TNIK::::5.7:C;MRCKA::::5.7:C;UFO::::5.7:C;PLK4::::5.7:C;FES::::5.7:C;MRCKB::::5.68:C;EPHA6::::5.68:C;EGFR:L858R-T790M:::5.66:C;EGFR:T790M:::5.64:C;TAOK3::::5.64:C;M3K10::::5.6:C;AURKA::::5.58:C;TGFR2::::5.54:C;M4K4::::5.51:C;FLT3:K663Q:::5.49:C;VRK2::::5.49:C;RET:V804L:::5.49:C;STK25::::5.47:C;MYLK2::::5.46:C;M3K7::::5.43:C;STK4::::5.42:C;ULK3::::5.34:C;FLT3::::5.32:C;FLT3:D835Y:::5.32:C;VGFR1::::5.3:C;PKN2::::5.3:C;IRAK4::::5.3:C;M3K13::::5.28:C;TAOK2::::5.27:C;NEK2::::5.19:C;WEE1::::5.15:C;FLT3:N841I:::5.15:C;BMR1A::::5.15:C;FLT3:D835H:::5.09:C;PUR1;HSP7C;BCR;NR4A3;STA5B:::inh::D|CP3A4:::inh:5.2:DC;FMO3:::sub::D;CP3A5:::sub::D;CP1B1:::sub::D;CP1A2:::sub::D;CP1A1:::sub::D|ABCG2:::inh::D;MDR1:::inh::D|
Lisdexamfetamine|ok_inv|TAAR1:::ago::D|CP2D6:::inh::D|S15A1:::sub::D|
Retapamulin|ok|RL3::STRP1:inh::D|CP3A4:::sub::D||
Eculizumab|ok_inv|CO5:::abo::D|||
Lapatinib|ok_inv|EGFR:G719C::ant:9.04:DC;EGFR:L861Q::ant:8.92:DC;ERBB2:::ant:8.8:DC;EGFR:G719S::ant:8.68:DC;EGFR:::ant:8.66:DC;EGFR:L858R::ant:8.55:DC;ERBB4::::7.6:C;TBA1A::RAT::7.27:C;P3C2B::::6.17:C;EGFR:T790M::ant:6.07:DC;PI4KB::::6.03:C;KCNH2::::6.:C;MP2K5::::5.96:C;RET::::5.9:C;AURKB::::5.7:C;STK10::::5.59:C;SLK::::5.48:C;RIPK2::::5.44:C;MP2K7::::5.36:C;ERBB3::::5.26:C;P3C2G::::5.12:C;PGFRB::::5.07:C|CP3A4:::inh:5.77:DC;CP2CJ:::sub::D;CP2C8:::inh::D;CP3A5:::sub::D|TAP1:::inh::D;MDR1:::inh::D|
Desonide|ok_inv|GCR:::ago::D|CP3A4:::sub_ind::D||
Sitagliptin|ok_inv|DPP4:::inh:8.46:DC;DPP8::::5.74:C;DPP9::::5.51:C;SEPR::::5.23:C|CP2C8:::sub::D;CP3A4:::sub::D|S22A8:::sub::D;MDR1:::sub::D|
Decitabine|ok_inv|DNMT1:::inh::D;DNA|DCK:::sub::D||
Posaconazole|ok_inv_vet|CP51::CANAL:ant::D|CP3A4:::inh:7.3:DC|MDR1:::inh::D|
Darunavir|ok|Pol_polyprotein::9HIV1:inh::D|CP3A4:::inh::D|MDR1:::inh::D;SO1B1:::inh::D|
Telbivudine|ok_inv|DNA;DPOL::HBVF1:::D|||
Sinecatechins|ok_inv_nutra||||
Paliperidone|ok|KCNH2::::6.:C;5HT7R;DRD1:::ant::D;5HT1A:::ant::D;ADA2C:::ago::D;ADA2B:::ant::D;ADA2A:::ant::D;5HT2C:::ant::D;DRD3:::ant::D;5HT1D:::ant::D;DRD4:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;HRH1:::ant::D;DRD2:::ant::D;5HT2A:::ant::D|CP3A5:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|
Sunitinib|ok_inv|PGFRB:::inh:10.12:DC;VGFR2:::inh:9.7:DC;KIT:V559D-V654A::inh:9.68:DC;FLT3:K663Q::inh:9.66:DC;KIT:V559D-T670I::inh:9.55:DC;KIT:::inh:9.43:DC;KIT:V559D::inh:9.39:DC;FLT3:::inh:9.39:DC;PGFRA:::inh:9.1:DC;ST17A::::9.:C;VGFR1:::inh:9.:DC;KIT:L576P::inh:8.89:DC;CSF1R:::inh:8.7:DC;FLT3:D835Y::inh:8.64:DC;FLT3:N841I::inh:8.62:DC;FLT3:D835H::inh:8.37:DC;BMP2K::::8.26:C;PHKG1::::8.26:C;RET:V804M:::8.24:C;PHKG2::::8.23:C;CHK2::::8.15:C;PGFRB::MOUSE::8.1:C;RET:V804L:::8.06:C;UFO::::8.05:C;VGFR3:::inh:8.05:DC;LCK::::8.05:C;JAK1::::8.05:C;AAK1::::7.96:C;FLT3:R834Q::inh:7.96:DC;RET::::7.92:C;KC1E::::7.89:C;ITK::::7.89:C;ULK2::::7.89:C;IRAK1::::7.85:C;KC1D::::7.82:C;MYLK4::::7.82:C;LRRK2::::7.82:C;M4K1::::7.8:C;PAK3::::7.8:C;STK33::::7.77:C;M3K19::::7.77:C;KS6A2::::7.77:C;KS6A5::::7.77:C;AAPK1::::7.72:C;STK10::::7.72:C;STK4::::7.72:C;RET:M918T:::7.72:C;CLK2::::7.7:C;GAK::::7.7:C;CLK1::::7.66:C;DAPK3::::7.66:C;ULK1::::7.64:C;MYLK::::7.64:C;MYLK::CHICK::7.64:C;MYLK3::::7.64:C;TNIK::::7.6:C;MERTK::::7.59:C;CLK4::::7.54:C;MINK1::::7.54:C;HIPK2::::7.51:C;M4K2::::7.48:C;RIOK1::::7.46:C;STK11::::7.42:C;PI42B::::7.41:C;M4K5::::7.39:C;HIPK3::::7.39:C;ULK3::::7.38:C;KIT:A829P::inh:7.37:DC;MP2K5::::7.34:C;NUAK1::::7.32:C;KS6B1::::7.32:C;TYRO3::::7.31:C;RIOK2::::7.31:C;MYLK2::::7.31:C;ABL1:T315I:::7.26:C;ALK::::7.26:C;KS6A3::::7.26:C;HIPK1::::7.26:C;STK3::::7.25:C;SLK::::7.25:C;M3K2::::7.24:C;SRPK3::::7.23:C;TTK::::7.2:C;STK24::::7.2:C;BLK::::7.19:C;IRAK4::::7.18:C;ABL1:H396P:::7.13:C;ABL1:Q252H:::7.12:C;LRRK2:G2019S:::7.12:C;CHK1::::7.11:C;KCC2A::::7.1:C;CSK21::::7.09:C;FAK2::::7.09:C;PKNB::MYCTU::7.06:C;AAPK2::::7.05:C;M3K7::::7.03:C;M3K13::::7.02:C;KS6A1::::7.02:C;KS6A4::::7.02:C;DLK1::::7.:C;NTRK1::::7.:C;KC1A::::7.:C;M3K12::::7.:C;KC1G2::::6.96:C;DCLK3::::6.96:C;ST17B::::6.96:C;MP2K2::::6.96:C;KIT:D816H::inh:6.96:DC;ULK3::MOUSE::6.96:C;DAPK1::::6.92:C;TBK1::::6.92:C;YES::::6.92:C;ABL1:M351T:::6.92:C;MP2K1::::6.89:C;CDK16::::6.89:C;M4K4::::6.85:C;GRK4::::6.85:C;STK39::::6.85:C;ROCK2::::6.85:C;ABL1:Y253F:::6.85:C;DAPK2::::6.82:C;NUAK2::::6.82:C;ABL1::::6.82:C;SRC::::6.82:C;HIPK4::::6.8:C;CSK22::::6.8:C;STK3::MOUSE::6.8:C;FGFR1::::6.77:C;EGFR::::6.76:C;GRK7::::6.74:C;M4K3::::6.74:C;E2AK4::::6.74:C;ABL1:E255K:::6.74:C;INSR::::6.74:C;SRPK2::::6.72:C;PLK4::::6.72:C;HCK::::6.72:C;DYR1A::::6.7:C;MAST1::::6.7:C;SBK1::::6.7:C;TAOK3::::6.68:C;AURKC::::6.66:C;M3K3::::6.66:C;SGK3::::6.66:C;KC1G3::::6.62:C;SRPK1::::6.6:C;STK16::::6.6:C;KCNH2::::6.6:C;FGR::::6.57:C;LYN::::6.57:C;CDK14::::6.57:C;KPCD3::::6.55:C;FGFR3::::6.54:C;RK::::6.54:C;STK25::::6.54:C;ANKK1::::6.51:C;MARK2::::6.51:C;KPCD1::::6.51:C;CDK7::::6.48:C;TLK2::::6.48:C;STK26::::6.47:C;MELK::::6.46:C;TYK2::::6.44:C;DCLK1::::6.43:C;RIPK1::::6.43:C;ABL1:F317L:::6.43:C;AURKB::::6.42:C;KPCD2::::6.42:C;KIT:D816V::inh:6.42:DC;PRP4::::6.41:C;PRP4B::::6.41:C;JAK2::::6.39:C;MARK3::::6.39:C;STK38::::6.39:C;KCC2D::::6.38:C;KKCC1::::6.38:C;INSRR::::6.37:C;KCC2G::::6.36:C;FAK1::::6.36:C;KCC1G::::6.36:C;LATS2::::6.34:C;ROCK1::::6.34:C;ICK::::6.33:C;EPHB1::::6.32:C;MUSK::::6.31:C;HUNK::::6.3:C;NEK2::::6.3:C;KCC1D::::6.29:C;FRK::::6.28:C;FYN::::6.28:C;IKKA::::6.28:C;OXSR1::::6.28:C;FGFR2::::6.28:C;KC1AL::::6.26:C;SRC::CHICK::6.26:C;BMPR2::::6.24:C;SIK2::::6.24:C;NTRK2::::6.23:C;ERN1::::6.22:C;IKKE::::6.21:C;LATS1::::6.2:C;PAK5::::6.19:C;SNRK::::6.19:C;DYRK2::::6.17:C;TNK1::::6.17:C;E2AK2::::6.17:C;PKN1::::6.15:C;MP2K4::::6.15:C;EPHA7::::6.15:C;TLK1::::6.13:C;EPHB6::::6.07:C;NIM1::::6.07:C;EGFR:L858R-T790M:::6.07:C;KCC4::::6.05:C;TAOK1::::6.05:C;ABL1:F317I:::6.05:C;KC1G1::::6.03:C;IRAK3::::6.03:C;EPHA6::::6.02:C;FES::::6.02:C;KCC1A::::6.01:C;ST38L::::6.01:C;ABL2::::6.:C;BRSK2::::5.96:C;CDKL2::::5.96:C;WEE1::::5.96:C;FER::::5.96:C;MARK1::::5.92:C;JAK3::::5.92:C;MET:M1250T:::5.92:C;EPHA5::::5.92:C;CDK17::::5.92:C;M3K15::::5.89:C;M3K11::::5.89:C;PKN2::::5.89:C;STK35::::5.89:C;DUSTY::::5.89:C;CDPK1::PLAF7::5.89:C;KCC2B::::5.85:C;FGFR3:G697C:::5.85:C;KKCC2::::5.82:C;AURKA::::5.77:C;CDK18::::5.77:C;MP2K3::::5.77:C;LTK::::5.74:C;SBK3::::5.72:C;DDR1::::5.7:C;MET::::5.7:C;CDK4::::5.7:C;EPHA3::::5.68:C;RIPK4::::5.68:C;FGFR4::::5.68:C;BTK::::5.68:C;EPHB4::::5.66:C;ACK1::::5.66:C;DYR1B::::5.64:C;PAK4::::5.64:C;PAK6::::5.62:C;PIM3::::5.62:C;KS6A6::::5.62:C;MK09::::5.62:C;BMR1B::::5.62:C;EGFR:T790M:::5.62:C;IGF1R::::5.59:C;DCLK2::::5.57:C;AKT2::::5.57:C;DDR2::::5.54:C;MYO3A::::5.51:C;SIK1::::5.49:C;M3K4::::5.48:C;M3K9::::5.47:C;BRSK1::::5.46:C;PDPK1::::5.46:C;MARK4::::5.44:C;RIOK3::::5.42:C;CTRO::::5.41:C;MKNK1::::5.41:C;TIE1::::5.41:C;NEK7::::5.39:C;KPCT::::5.37:C;MK10::::5.37:C;MYO3B::::5.35:C;PTK6::::5.34:C;PLK2::::5.33:C;MET:Y1235D:::5.33:C;PIM2::::5.3:C;NTRK3::::5.29:C;MP2K6::::5.28:C;PI51A::::5.27:C;MKNK2::::5.24:C;ACES::::5.23:C;KPCA::::5.22:C;MEN1::::5.2:C;TSSK1::::5.2:C;EGFR:G719C:::5.17:C;CDK5::::5.16:C;LMNA::::5.15:C;MATK::::5.11:C;TNKS2::::5.05:C;MK07::::5.:C|CP3A4:::inh::D;CP3A7:::sub::D;CP3A5:::sub::D|ABCG2:::inh::D;MRP2:::inh::D;MDR1:::inh::D;MRP4:::inh::D|
Panitumumab|ok_inv|EGFR:::sup::D|||
Ranibizumab|ok|VEGFA|||
Idursulfase|ok|Dermatan_sulfate;Heparan_sulfate;PLIN3|||
Alglucosidase_alfa|ok|MPRD:::bin::D;Glycogen:::cli::D|||
Varenicline|ok_inv|ACHA4::RAT::10.3:C;ACHB2:::pag:10.22:DC;ACHA2::RAT::9.66:C;ACHA3::RAT::8.72:C;ACHA7::RAT::7.49:C;ACHB3::RAT::7.34:C;ACHB4::::7.13:C;ACHA7:::ago:6.9:DC;ACHA::::5.09:C;ACHA6:::pag::D;ACHA3:::pag::D;ACHA4:::pag::D||S22A2:::inh::D|
Arformoterol|ok_inv|ADRB2::CAVPO::9.9:C;ADRB2:::ago:9.5:DC;ADRB3::::7.6:C;ADRB1::::7.4:C|CP2C9:::sub::D;CP2A6:::sub::D;CP2CJ:::sub::D;CP2D6:::sub::D||
Hydralazine|ok|ACM1::RAT::7.55:C;TPO::::7.4:C;PERM::::6.05:C;CP1A2::::6.:C;P53::::5.8:C;KPYK::LEIME::5.7:C;RAB9A::::5.64:C;NPC1::::5.59:C;LMNA::::5.5:C;LOX15::RABIT::5.44:C;LUCI::PHOPY::5.4:C;SMN::::5.4:C;FFP::BACIU::5.3:C;AL1A1::::5.3:C;KPYM::::5.1:C;HIF1A:::ind::D;P4HA1:::inh::D;AOC3:::inh::D|CP3A4:::inh:5.4:DC||ALBU:::bin::D
Exenatide|ok_inv|GLP1R:::ago:10.:DC;GLP1R::RAT::9.85:C|DPP4:::sub::D||ALBU
Mecasermin|ok_inv|IGF1R:::ago::D;IBP3;INSR;MPRI|||IBP3:::car::D;ALS:::car::D;IBP1:::car::D;IBP2:::car::D;IBP4:::car::D;IBP5:::car::D;IBP6:::car::D
Pramlintide|ok_inv|CALCR:::ago::D;RAMP1:::ago::D;RAMP2:::ago::D;RAMP3:::ago::D|||
Galsulfase|ok_inv|Dermatan_sulfate;PLIN3|||
Nelarabine|ok_inv|DPOLA:::inh::D;DNA:::destbz::D|DGUOK:::sub::D;DCK:::sub::D;ADA:::sub::D||
Abatacept|ok|CD80:::ant::D;CD86:::ant::D|||
Carbetocin|ok_inv|OXYR:::ago:9.15:DC;V1AR::::7.39:C;V2R::::6.77:C|||
Lumiracoxib|ok_inv|PGH1:::inh:8.15:DC;PGH2:::inh:8.15:DC;PGH2::MOUSE::7.4:C|CP1A2:::sub::D;UD19:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D||
Tetracosactide|ok|MC4R::::9.19:C;ACTHR:::ant::D|||
Corticotropin|ok_inv_vet|ACTHR:::ago::D;CRF:::ago::D|3BHS2:::ind::D;CP27B:::ind::D;CP24A:::ind::D;CP3A4:::sub_ind::D||
Fenoterol|ok_inv|ADRB2::CAVPO::7.74:C;ADRB2:::ago:7.:DC;ADRB3:::ago::D;ADRB1:::ago::D|||
Glisoxepide|inv|KCNJ8:::inh::D|CP2C9:::sub::D||
Pirbuterol|ok|ADRB2:::ago::D;ADRB1:::ago::D|||
Bismuth_subsalicylate|ok_vet||||ALBU:::bin::D;TRFE
Bevantolol|exp|ADRB1:::ant::D;ADRB2:::ant::D;ADA1A:::ant::D|CP2D6:::sub::D||
Glucosamine|ok_inv|TNFA;MMP9:::ant::D;NFKB2:::ant::D;IFNG;CHIS::BACCI:::D|||
Practolol|ok|ADRB2::CANLF::6.73:C;ADRB1:::ant:6.6:DC;ADRB1::RAT::6.47:C;ADRB2::CAVPO::5.8:C|CP2D6:::sub::D||
Sulfacytine|ok|DHPS::ECOLI:inh::D|||
Sulfadoxine|ok_inv|DRTS::PLAFK:inh::D;Dihydropteroate_synthetase::PLAFA:::D|||
Rolitetracycline|ok|16S_ribosomal_RNA::Gut_flora:inh::D;RS9::ECOLI:inh::D|||
Oxtriphylline|ok|PDE3A:::inh::D;PDE4A:::inh::D;AA2AR:::ant::D;AA1R:::ant::D;HDAC2:::act::D|CP1A2:::sub::D|S22A7:::inh::D|
Insulin_aspart|ok|INSR:::ago::D;IGF1R|CP1A2:::ind::D||
Insulin_detemir|ok|INSR:::ago::D;IGF1R|CP1A2:::ind::D||ALBU
Insulin_glulisine|ok|INSR:::ago::D;IGF1R|CP1A2:::ind::D||
Fosamprenavir|ok|Pol_polyprotein::9HIV1:inh::D|CP3A4:::inh::D||
Fosphenytoin|ok_inv|SCN5A:::inh::D|UD19:::inh::D;UD16:::inh::D;CP1A2:::ind::D;CP2B6:::ind::D;CP3A4:::sub_ind::D;CP2CJ:::sub::D;CP2C9:::sub_ind::D||THBG:::sub::D;ALBU
Josamycin|inv|RL4::HAEIN:inh::D|||
Kava|ok_inv_nutra||||
St_John_s_Wort|ok_inv_nutra||CP3A4:::sub_ind::D;CP2D6:::inh::D;CP2CJ:::sub_ind::D|MDR1:::ind::D|
Polythiazide|ok|S12A3:::inh::D|||
Quinethazone|ok|S12A3:::inh::D;S12A2:::inh::D;S12A1:::inh::D;CAH2:::inh::D;CAH1:::inh::D|||
Cefamandole|ok_exp|Penicillin_binding_protein_2::BACFG:inh::D||S22A6:::inh:7.52:DC;S22A8:::inh:7.34:DC;S22AB:::inh:5.94:DC;S22A7:::inh::D|
Cefazolin|ok|LMNA::::6.05:C;IL2:::inh::D;IL15:::inh::D;PON1:::inh::D;FTSI::ECOLI:inh::D;MRDA::ECOLI:inh::D;PBPC::ECOLI:inh::D;PBPB::ECOLI:inh::D;PBPA::ECOLI:inh::D|TPMT:::sub::D|S22A6:::inh:6.74:DC;S22A8:::inh:6.26:DC;S22AB:::inh:5.76:DC;MRP4:::sub::D|ALBU
Cefonicid|ok_inv|MRDA::ECOLI:inh::D;DACB::ECOLI:inh::D;PBPB::ECOLI:inh::D;FTSI::ECOLI:inh::D;PBPA::ECOLI:inh::D|||ALBU
Cefoperazone|ok_inv|DACB::ECOLI:inh::D;DACA::ECOLI:inh::D;PBPA::ECOLI:inh::D;DACC::ECOLI:inh::D;Penicillin_binding_protein_1B::PSEAI:inh::D;PBPA::PSEAE:inh::D;MRDA::ECOLI:inh::D;PBPB::ECOLI:inh::D;FTSI::ECOLI:inh::D||S22A6:::inh:6.68:DC;S22A8:::inh:5.72:DC;S22AB:::inh:5.55:DC;S22A7:::inh::D|ALBU
Cefotetan|ok|LMBL1::::5.1:C;PBP3::STREE:inh::D|||ALBU
Cefoxitin|ok|PBP2::STRR6:inh::D;PBPA::STRR6:inh::D;PBP2A::STRR6:inh::D;PBP1B::STRR6:inh::D;PBP3::STREE:inh::D;FTSI::ECOLI:inh::D;PBPB::ECOLI:inh::D;PBPA::ECOLI:inh::D;DACB::ECOLI:inh::D;PBP7::ECOLI:inh::D;DACA::ECOLI:inh::D;DACC::ECOLI:inh::D|BLAC::BACLI:sub::D||
Ceftizoxime|ok_inv|MecA::STAAU:inh::D;PBPA::ECOLI:inh::D;PBPB::ECOLI:inh::D;FTSI::ECOLI:inh::D||S15A1:::sub::D;S22A6:::sub::D;S22A8:::inh::D|
Cefradine|ok|PBPA::ECOLI:inh::D|CP3A4:::ind::D|S15A1:::inh:5.01:DC;S47A1:::sub::D;S22A6:::inh::D;S15A2:::inh::D;S22A5:::inh::D|
Metocurine|ok|ACM2:::ant::D;ACHA2:::ant::D|||
Pancuronium|ok|MTOR::::6.68:C;ACM3:::ant::D;ACM2:::ant::D;ACHA2:::ant::D|CHLE:::inh::D|S22A2;S22A1:::sub::D|
Pipecuronium|ok|ACHA2:::ant::D;ACM2:::ant::D;ACM3:::ant::D|CHLE:::inh::D||
Vecuronium|ok_inv|ACHA2:::ant::D||MDR1:::sub::D|
Cilazapril|ok|ACE:::inh::D||S15A2:::sub::D;S15A1:::sub::D;MDR1:::inh::D|
Tolevamer|ok_inv|Potassium:::bin::D|||
Potassium_cation|ok_inv|AT1A1|||
Quinidine_barbiturate|ok|GBRA1:::pot::D;GBRA2:::pot::D;SCN5A:::inh::D;KCNK1:::inh::D;GRIA2:::ant::D|||
Spirapril|ok|ACE::RAT::7.17:C;ACE:::inh::D||S15A2:::sub::D;S15A1:::sub::D|
Tasosartan|exp|AGTRB::RAT::8.92:C;AGTR1:::ant:8.4:DC;AGTR2:::ant::D|CP3A4:::sub::D||
Amobarbital|ok_ill|GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|||
Aprobarbital|exp_ill|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA4:::pot::D;GBRA5:::pot::D;GBRA6:::pot::D;ACHA4:::ant::D;ACHA7:::ant::D;GRIA2:::ant::D;GRIK2:::ant::D|CP3A4:::ind::D||
Butobarbital|ok_ill|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA4:::pot::D;GBRA5:::pot::D;GBRA6:::pot::D;ACHA4:::ant::D;ACHA7:::ant::D;GRIA2:::ant::D;GRIK2:::ant::D|||
Heptabarbital|exp|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA4:::pot::D;GBRA5:::pot::D;GBRA6:::pot::D;ACHA4:::ant::D;ACHA7:::ant::D;GRIA2:::ant::D;GRIK2:::ant::D|||
Hexobarbital|exp|MEN1::::5.55:C;GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|PGH1:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D||
Mestranol|ok|ESR1:::ago:8.28:DC;SC6A4::::7.66:C;LMNA::::5.9:C;SC6A2::::5.86:C;ANDR::RAT::5.15:C;RORG::MOUSE::5.15:C|CP2C8:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D||
Penbutolol|ok_inv|5HT1A::RAT::8.62:C;5HT1B:::ant::D;5HT1A:::ant::D;ADRB2:::ant_pago::D;ADRB1:::ant_pago::D|CP2D6:::sub::D||A1AG1
Iohexol|ok||||
Ephedrine|ok|ACES;VMAT2:::inh::D;ADA1A;SC6A2:::ANT::D|CHLE:::sub::D||
Mephentermine|ok|LMNA::::8.49:C;CP2D6::::5.:C;ADRB1,ADRB2,ADRB3:::ago::D;ADA1A,ADA1B,ADA1D,ADA2A,ADA2B,ADA2C:::ago::D|||
Procaterol|ok_inv|TSHR::::7.9:C;ADRB2:::ago:7.48:DC|||
Rasagiline|ok|AOFA::RAT::9.:C;AOFB:::inh:8.4:DC;AOFB::RAT::8.36:C;AOFA::::6.39:C;BCL2:::act::D|CP1A2:::sub::D||
Quinupristin|ok|23S_ribosomal_RNA::Gut_flora:inh::D;RL10::SHIFL:inh::D;RL22::ECO57:inh::D|CP3A4:::inh::D||
Aluminium|ok_inv|TRFE;AT1A1:::bin::D;KLK1:::inh::D;A4|||ALBU
Calcium|ok_nutra|CAC1C:::lig::D;AT2C1:::ago::D;TNNC2:::ago::D;TNNC1:::ago::D;SPTB2:::ago::D;S100B;ICAL;COMP;CALM1;AOC1;S10AD;PPB1;S10A8;S10A9;S10A2;CERU;BMP4;MGP;PCD19;PDCD6|||
Magnesium_oxide|ok||||
Magnesium_cation|ok_nutra|AT1A1|||
Cortisone_acetate|ok_inv|GCR:::ago:5.75:DC;ACM1::RAT::5.:C|CP3A5:::ind::D;CP3A4:::sub_ind::D||
Ginkgo_biloba|ok_inv_nutra|SC6A2:::inh::D;PA2GA:::inh::D;GLRA1:::ant::D;GBRA1:::neg::D;GBRB2:::neg::D;GBRG2:::neg::D|CP2C9:::inh::D;CP3A4:::inh::D||
Glymidine|ok_inv|KCNJ1;ABCC8:::ind::D|||
Paramethasone|exp|GCR:::ago::D|CP3A5:::ind::D;CP3A4:::duo::D||CBG:::bin::D
Mibefradil|inv_out|CAC1H:::inh:7.49:DC;CAC1I:::inh:6.9:DC;CAC1C:::inh:6.81:DC;KCNH2::::6.72:C;CAC1G:::inh:6.7:DC;CAC1B::::6.38:C;SCN1A::::6.01:C;CAC1C::RAT::5.96:C;CP2CJ::::5.88:C;CP2J2::::5.67:C;TAU::::5.55:C;MDR1A::MOUSE::5.13:C;MDR1B::MOUSE::5.:C;CACB4:::inh::D;CACB3:::inh::D;CACB2:::inh::D;CACB1:::inh::D;CAC1S:::inh::D;CAC1F:::inh::D;CAC1D:::inh::D|CP2D6:::inh:7.2:DC;CP3A4:::inh:6.89:DC;C11B2:::inh::D;C11B1:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP1A2:::inh::D|MDR1:::inh:5.92:DC|
Sodium_bicarbonate|ok|Hydrogen_ions::UNK:neu::D||S4A10:::sub::D;S4A5:::sub::D;S4A8:::sub::D;S4A7:::sub::D;S4A4:::sub::D|
Yohimbine|ok_inv_vet|ADA2A:::ant:9.4:DC;ADA2C:::ant:9.3:DC;ADA2B::MOUSE::9.22:C;ADA2C::RAT::9.22:C;ADA1B::::8.96:C;ADA1D::::8.8:C;ADA2B::RAT::8.7:C;ADA2B:::ant:8.7:DC;ADA1A::BOVIN::8.44:C;ADA2A::PIG::8.36:C;ADA1B::RAT::8.14:C;CAC1C::RAT::7.35:C;5HT2B:::ant:7.33:DC;ADA2A::BOVIN::7.31:C;ADA1D::RAT::7.28:C;5HT1A::RAT::7.14:C;AA3R::::7.02:C;ADA1A::::6.83:C;ADA1A::RAT::6.3:C;DRD2:::ant:6.16:DC;5HT6R::::6.11:C;DRD2::RAT::5.95:C;5HT2A::RAT::5.79:C;DRD5::RAT::5.7:C;DRD3::RAT::5.61:C;KCNJ1,KCJ10,KCJ11,KCJ12,KCJ14,KCJ15,KCNJ8:::inh::D;5HT2C:::ant::D;5HT2A:::ant::D;DRD3:::ant::D;5HT1D:::ant::D;5HT1B:::ant::D;5HT1A:::pag::D|CP2D6:::sub:8.08:DC;CP3A4:::sub::D||
Bezafibrate|ok_inv|PPARG:::ago:5.98:DC;PPARA:::ago:5.15:DC;RXRG:::ago::D;RXRB:::ago::D;RXRA:::ago::D;NR1I2:::pag::D;PPARD:::ago::D|CP3A4:::sub::D;CP2C8:::inh::D;CP1A1:::ind::D|SO1B1:::inh::D|
Colchicine|ok|MITF::::7.25:C;TBB5:::inh::D|CP2E1:::ind::D;CP2C8:::inh::D;CP2B6:::inh::D;CP3A4:::inh::D|MDR1:::sub_ind::D|ALBU:::bin::D
Drospirenone|ok|GCR:::bin::D;ANDR:::ant::D;MCR:::ant::D;PRGR:::ago::D|CP3A4:::sub::D;PON1:::sub::D;PGH2:::duo::D||
Digitoxin|ok_inv|AT1A1:::inh:8.1:DC;AT1A1::CANLF::8.1:C;P53::::7.5:C;LMNA::::6.15:C;STAT3::::6.15:C;RORG::MOUSE::5.95:C;CYSP::TRYCR::5.7:C;TAU::::5.15:C|CP11A:::inh::D;CP3A4:::sub::D|SO4C1:::inh:6.92:DC;MDR1:::sub::D;SO1A2:::inh::D|ALBU
Salsalate|ok|PGH1:::inh::D;PGH2:::inh::D|||
Neostigmine|ok_vet|ACES::TETCF::8.34:C;ACES:::inh:5.62:DC;LMNA::::5.3:C;ACM1::RAT::5.25:C|CHLE:::inh::D||
Choline_magnesium_trisalicylate|ok|PGH1:::inh::D;PGH2:::inh::D|||
Methotrimeprazine|ok_inv|PDR5::YEAST::5.02:C;ADA2C:::ant::D;ADA2B:::ant::D;ADA2A:::ant::D;ADA1D:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;HRH1:::ant::D;5HT2C:::ant::D;5HT2A:::ant::D;DRD4:::ant::D;DRD3:::ant::D;DRD5:::ant::D;DRD1:::ant::D;DRD2:::ant::D|CP2E1:::inh::D;CP2D6:::inh::D||
Ginseng|ok_inv_nutra|IL6:::ant::D;PGH2:::inh::D;AHR:::ago::D|||
Temafloxacin|out|PARC::HAEIN:inh::D;GYRA::HAEIN:inh::D|CP1A2:::inh::D||
Danazol|ok|ANDR::RAT::8.1:C;CP2J2::::7.92:C;CP2C9::::6.52:C;GCR::::5.71:C;CP2C8::::5.71:C;5HT2A::::5.6:C;CP2D6::::5.56:C;ADA2C::::5.46:C;ACM3::::5.42:C;ESR1:::ago:5.29:DC;SC6A3::::5.26:C;SC6A2::::5.25:C;OPRM::::5.24:C;OPRK::::5.21:C;AA3R::::5.2:C;ADA2A::::5.16:C;SC6A4::::5.09:C;NK2R::::5.05:C;DRD3::::5.01:C;CCL2:::inh::D;GNRR2:::neg::D;GNRHR:::neg::D;PRGR:::ago::D;ANDR:::ago::D|CP3A4:::inh::D;CP19A:::inh::D||SHBG:::ant:8.2:DC
Clenbuterol|ok_inv_vet|ADRB2::CAVPO::7.89:C;ADRB2:::ago:7.8:DC;ADRB2::BOVIN::7.44:C;ADRB1:::ago:7.16:DC;5HT1A::RAT::5.82:C;TNFA;NGF:::sti::D;ADRB3:::ago::D|CP1A1:::sub::D||
Bambuterol|inv|CP2D6::::5.7:C;AMPC::ECOLI::5.3:C;ADRB2:::ago::D|CHLE:::inh::D||
Tiotropium|ok|ACM5;ACM4;ACM2:::ant::D;ACM1:::ant::D;ACM3:::ant::D|CP3A4:::sub::D;CP2D6:::sub::D|S22A4:::sub::D;S22A5:::sub::D|
Ciclesonide|ok_inv|GCR:::ago::D|EST1:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D||CBG:::bin::D
Pranlukast|inv|CLTR1:::ant:10.36:DC;CLTR1::CAVPO::9.1:C;CLTR2::::5.44:C;GPR17::::5.39:C;CYSP::TRYCR::5.15:C;MUC2;NFKB1;ECP;IL5:::ant::D;TNFA|CP2C9:::inh::D;CP3A4:::sub::D|MRP2:::inh::D|
Theobromine|inv|ACM1::RAT::7.95:C;PDE4B:::inh::D;AA2AR:::ant::D;AA1R:::ant::D|CP2E1:::sub::D;CP1A2:::sub::D||
Cefepime|ok_inv|Penicillin_binding_protein_2::PSEAI:inh::D;Cell_division_protein::PSEAI:inh::D;FTSI::ECOLI:inh::D;MRDA::ECOLI:inh::D||S15A2:::inh::D;S15A1:::inh::D;S22A5:::inh::D|
Cefacetrile|exp_vet|PBPA::ECOLI:inh::D;PBPB::ECOLI:inh::D||S22A6:::inh::D;S22A8:::inh::D|
Ceftibuten|ok_inv|MRDA::ECOLI:inh::D;PBPB::ECOLI:inh::D;PBPA::ECOLI:inh::D;FTSI::ECOLI:inh::D||S22A8:::inh::D;S22A6:::sub::D;S15A2:::inh::D;S15A1:::inh::D|
Cefpodoxime|ok_vet|FTSI::ECOLI:inh::D|||
Acenocoumarol|ok_inv|VKOR1:::inh::D|CP3A4:::sub::D;CP2CJ:::sub::D;CP1A2:::sub::D;CP2C9:::sub::D|MDR1:::sub::D|A1AG1;ALBU
Antrafenine|ok|PGH1:::inh::D;PGH2:::inh::D|||
Testosterone_propionate|ok_inv_vet_out|ANDR:::ago:9.6:DC;ANDR::MOUSE::8.55:C;LMNA::::8.1:C;CP17A::::7.25:C;ANDR::RAT::5.72:C;CP2CJ::::5.:C|CP3A4:::sub:5.9:DC;S5A1,S5A2,PORED:::sub::D;UD11:::ind::D;COMT:::inh::D|MDR1:::sub::D|ALBU:::sub::D;SHBG:::sub::D
Paromomycin|ok_inv|16S_ribosomal_RNA::Gut_flora:inh::D;RS10::THET8:inh::D|||
Nitroxoline|exp|MAP2:::inh:7.26:DC;RORG::MOUSE::6.55:C;LMNA::::6.05:C;HS90A::::6.:C;PGH2::::6.:C;KDM4E::::5.55:C;HD::::5.45:C;DNAB::MYCTU::5.18:C;TAU::::5.05:C;Manganese_cation:::chel::D;Magnesium_cation:::chel::D|||
Stepronin|exp||||
Aminophenazone|ok_out|LMNA::::7.2:C;TSHR::::5.1:C|CP1A2:::sub:5.:DC;CP17A:::sub::D;CP2CI:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::inh::D|S22A6:::inh::D|
Alizapride|inv|DRD2::RAT::6.7:C;DRD2:::ant::D|||
Ajmaline|ok_exp|SCN5A:::inh::D|||A1AG1
Amrinone|ok|LMNA::::6.5:C;HD::::6.3:C;KDM4E::::5.95:C;HCD2::::5.9:C;AGAL::::5.9:C;TAU::::5.85:C;CP3A4::::5.5:C;HIF1A::::5.4:C;PDE4A::::5.32:C;CP2CJ::::5.3:C;FFP::BACIU::5.25:C;MEN1::::5.2:C;PDE3B:::inh::D;TNFA:::inh::D;PDE4B:::inh::D;PDE3A:::inh::D|||
Oxybenzone|ok_inv|CP2CJ::::6.4:C;CP1A2::::5.8:C;LIPS::RAT::5.49:C;PGDH::::5.05:C;ESR2;ESR1;ANDR:::ant::D;PRGR:::ant::D|||
Aprindine|exp|CALM1:::inh::D;SCN5A:::inh::D|CP2D6:::sub::D||A1AG1
Almitrine|ok|AT1A1:::bin::D|||
Allylestrenol|exp|ESR1:::ago::D;PRGR:::ago::D|||
Cholestyramine|ok_inv|Bile_acids:::bin::D|||
Antipyrine|ok_inv|PGH1:::inh::D;PGH2:::inh::D|CP2E1:::sub::D;CP2D6:::sub::D;CP2CI:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;CP3A4:::sub::D;CP2CJ:::sub::D;CP1A2:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D|S22A6:::inh::D|
Alfacalcidol|ok_nutra|SC6A2::::6.:C;RXRA;CP27B;VDR:::ago::D|||VTDB:::sub::D
Glutethimide|ok_ill|GABAR:::aga::D;GBRA1:::ago::D|CP11A:::inh::D||
Phenazopyridine|ok|Group_A_nerve_fibers::Rat:inh::D;SCN1A:::inh::D|||
gamma_Hydroxybutyric_acid|ok_ill_inv|S52A2:::ago::D;GBRB1:::ago::D||MOT2:::inh::D;MOT1:::inh::D;MOT4:::sub::D|
Diamorphine|ok_ill_inv|OPRM:::ago::D;OPRK:::ago::D;OPRD:::ago::D;EST1|||THBG:::ind::D
Bezitramide|exp_ill_out||||
Fencamfamin|exp_ill_out|SC6A3:::inh::D|||
Ethylmorphine|exp_ill|OPRM:::ago::D|CP3A4:::sub::D;CP2B6:::sub::D;NCPR:::ind::D;CP2D6:::sub::D||
Fenethylline|exp||CP1A2:::sub::D||
Barbital|ill|GRIK2:::ant::D;GRIA2:::ant::D;ACHA7:::ant::D;ACHA4:::ant::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2CJ:::sub_ind::D;CP3A4:::ind::D||
Cathine|exp_ill|HIF1A::::5.2:C;LMNA::::5.1:C|||
Camazepam|exp_ill||||
Ethylestrenol|out|ANDR::RAT::7.74:C;SC6A4::::7.37:C;ACM2::::6.98:C;ESR1::::6.49:C;CP2CJ::::5.89:C;SC6A2::::5.68:C;ACES::::5.19:C|||
Dichloralphenazone|ok_ill||||
Difenoxin|ok_ill||||
Dextromoramide|exp_ill||||
Chlorhexadol|exp_ill||||
Acetyldihydrocodeine|exp_ill||||
Flunitrazepam|ok_ill|GBRG2:::ago:8.96:DC;GBRA1:::ago:8.85:DC;GBRP::RAT::8.82:C;GBRA5:::pot:8.52:DC;GBRB3:::ago::D;GBRA3:::pot::D;GBRA6:::pot::D;GBRA4:::ago::D;GBRA2:::pot::D;TSPO:::ago::D|UD13:::inh::D;UD11:::inh::D;CP2E1:::inh::D;CP3A4:::sub::D;CP2C9:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;UD2B7:::inh::D;CP2CJ:::sub::D||
Ethyl_loflazepate|exp_ill||||
Dihydrocodeine|ok_ill||CP3A4:::sub::D;CP2D6:::sub::D||
Cloxazolam|exp|AK1C3::::5.82:C|||
Bromazepam|ok_ill_inv|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA4:::pot::D;GBRA5:::pot::D;GBRA6:::pot::D;GBRB1:::pot::D;GBRB2:::pot::D;GBRB3:::pot::D;GBRG1:::pot::D;GBRG2:::pot::D;GBRG3:::pot::D;GBRD:::pot::D;GBRE:::pot::D;GBRP:::pot::D;GBRR1:::pot::D;GBRR2:::pot::D;GBRR3:::pot::D;GBRT:::pot::D|CP1A2:::sub::D;CP2CJ:::sub::D;CP2E1:::inh::D||
Clotiazepam|ok_ill|GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRA5:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP3A4:::sub::D;CP2CJ:::sub::D;CP2CI:::sub::D;CP2B6:::sub::D||
Chloral_hydrate|ok_ill_inv_vet||||
Fludiazepam|exp_ill|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA5:::pot::D;GBRG1:::pot::D;GBRG2:::pot::D;GBRG3:::pot::D;GBRB1:::pot::D;GBRB2:::pot::D;GBRB3:::pot::D;GBRD:::pot::D;GBRE:::pot::D;GBRP:::pot::D;GBRR1:::pot::D;GBRR2:::pot::D;GBRR3:::pot::D|||
Attapulgite|ok_vet||||
Kaolin|ok||||
Dextroamphetamine|ok_ill|TAAR1::MOUSE::8.7:C;SC6A2:::neg:8.15:DC;SC6A3::RAT::7.61:C;TAAR1::RAT::7.25:C;TAAR1:::ago:6.85:DC;TAAR1::MACMU::6.:C;SC6A4::::5.75:C;SC6A4::RAT::5.75:C;5HT3A::RAT::5.35:C;ADA1B:::ant::D;ADA1A;VMAT2:::ind::D|AMO::ECOLI:sub::D;CP2D6:::sub::D|SC6A3::::7.61:DC|
Metamfetamine|ok_ill|TAAR1::MOUSE::7.15:C;TAAR1::RAT::6.88:C;TAAR1:::ago:5.89:DC;VMAT2::RAT::5.61:C;TAAR1::MACMU::5.28:C;SGMR1::::5.08:C;AOFB:::inh::D;AOFA:::inh::D;ADA2C:::ago::D;ADA2B:::ago::D;ADA2A:::ago::D;VMAT1:::inh::D;VMAT2:::inh::D;SC6A2:::neg::D;SC6A4:::neg::D;SC6A3:::neg::D|CP2D6:::sub::D|S22A5:::inh::D;S22A3:::inh::D|
Metrizamide|exp|AMPC::ECOLI::5.2:C|||
Phendimetrazine|ok_ill|ADA1B:::ago::D;SC6A2:::neg::D;ADA1A:::ago::D|||
Oxprenolol|ok|5HT1A::RAT::7.03:C;ADRB3;ADRB2:::ant::D;ADRB1:::ant::D|CP2D6:::inh::D|S22A2:::inh::D|
Sulfamerazine|ok_vet|DHPS::ECOLI:inh::D|||ALBU
Sulfamethazine|ok_inv_vet|DHPS::ECOLI:inh::D|NAT::MYCTU:sub::D||ALBU
Liotrix|ok|THA:::ago::D;THB:::ago::D|CP2C8:::inh::D;CP3A4:::sub::D|SO1A2:::sub::D;SO1B1:::sub::D;SO1B3:::sub::D;SO4C1:::sub::D;NTCP:::sub::D;SO1C1:::inh::D;SO4A1:::inh::D;S22A8:::inh::D;MOT8:::inh::D;MOT10:::inh::D;MDR1:::ind::D|TTHY;THBG:::sub::D;ALBU
Thyroglobulin|ok_out||||
Ursodeoxycholic_acid|ok_inv|CISD1::::5.95:C;GPBAR::::5.62:C;NR1H4;AK1C2:::ind::D|CP2E1:::duo::D|NTCP:::inh:5.44:DC;NTCP2:::inh::D;MRP4:::inh::D;MRP2:::ind::D;SO1A2:::duo::D;ABCBB:::duo::D|
Ketazolam|ok|TSPO:::ago::D;GBRA1:::pot::D;GBRB1:::pot::D;GBRG1:::pot::D;GBRD:::pot::D;GBRE:::pot::D|CP3A4:::inh::D|MDR1:::sub::D|ALBU
Prazepam|ok_ill|GABAR:::aga::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRA5:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP3A4:::sub::D||
Quazepam|ok_ill|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA5:::pot::D;GBRG1:::pot::D;GBRG2:::pot::D;GBRG3:::pot::D;GBRB1:::pot::D;GBRB3:::pot::D;GBRD:::pot::D;GBRE:::pot::D;GBRP:::pot::D;GBRR1:::pot::D;GBRR2:::pot::D;GBRR3:::pot::D;GABAR:::aga::D|CP2CJ:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D;CP2B6:::inh::D||
Everolimus|ok|MTOR:::inh::D|CP2D6:::inh::D;CP3A4:::sub::D|SO1A2:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D|
Solifenacin|ok|ACM1::RAT::8.:C;ACM3::RAT::8.:C;ACM2::RAT::6.92:C;KCNH2::::6.6:C;CAC1C::::5.37:C;SCN5A::::5.2:C;ACM5:::ant::D;ACM4:::ant::D;ACM2:::ant::D;ACM1:::ant::D;ACM3:::ant::D|CP2D6:::sub::D;CP1A1:::sub::D;CP3A4:::sub::D||A1AG1,A1AG2:::bin::D
Iron|ok|TFR1;EGLN1;HDAC8:::cof::D;AHSP;HBA;FRDA;FRIH;FEN1;NEIL1;NEIL2;DPOLB;CERU;TRFE|||
Zinc|ok_inv|BKRB1;MGMT;ALDOA;EF1A1;ENOA;G3PT;NDKA;PDIA1;PDIA3;PRDX1;SERB;TPIS;EFTU;ESR1:::cof::D;IL3;MT2;CCS;HDAC1:::cof::D;HDAC4:::cof::D;3MG;SEMG1;SODC;HDAC8:::cof::D;SIVA;GLRA1;MDM2;INS;UTRO;ACY2:::cof::D;S10A8;S10A9;MMP9;P73:::cof::D;S10A2;P53;MT3;PDCD6;DAND5:::cof::D;MT1A;A1BG;A2MG;ANGT;FETUA;SAMP;APOA1;APOA2;APOA4;APOBR;APOE;APOL1;C1QB;C1QC;C1R;C1S;CO3;CO4B;C4BPA;C4BPB;CO5;BRCC3;CO8A;CO8B;CO8G;CFAB;CFAH;CFAI;CLUS;CERU;CBPN;CPN2;DCD;DESP;FA12;F13B;THRB;FCN3;FIBA;FINC;GELS;HBA;HBB;HPTR;HORN;ALS;IGHA1;IGHM;KV117;KV320;LV321;ITIH1;ITIH2;ITIH3;ITIH4;IGJ;PLAK;KLKB1;KNG1;K2C1;K1C10;K1C14;K1C16;K22E;K2C5;K2C6A;K1C9;A1AG2;PGRP2;PON1;PZP;S10A7;SEPP1;A1AT;AACT;KAIN;CBG;HEP2;SHBG;TRFE;TTHY;VTNC;APLP1:::cof::D;APLP2:::cof::D;A4:::cof::D;PARP1|CAH1:::sub::D||
Cinolazepam|exp|GBRA1:::pot::D;GBRA2:::pot::D;GBRA3:::pot::D;GBRA5:::pot::D;GBRG1:::pot::D;GBRG2:::pot::D;GBRG3:::pot::D;GBRB1:::pot::D;GBRB2:::pot::D;GBRB3:::pot::D;GBRD:::pot::D;GBRE:::pot::D;GBRP:::pot::D;GBRR1:::pot::D;GBRR2:::pot::D;GBRR3:::pot::D|||
Nitrazepam|ok|GBRA2::BOVIN::7.42:C;LMNA::::5.45:C;SCN1A;GBRT:::pot::D;GBRR3:::pot::D;GBRR2:::pot::D;GBRR1:::pot::D;GBRP:::pot::D;GBRE:::pot::D;GBRD:::pot::D;GBRG3:::pot::D;GBRG2:::pot::D;GBRG1:::pot::D;GBRB3:::pot::D;GBRB2:::pot::D;GBRB1:::pot::D;GBRA6:::pot::D;GBRA5:::pot::D;GBRA4:::pot::D;GBRA3:::pot::D;GBRA2:::pot::D;GBRA1:::pot::D|CP2E1:::inh::D;CP3A4:::sub::D||
Cilastatin|ok_inv|DPEP1::PIG::6.96:C;DPEP1:::inh::D||S22A8:::inh::D;S22A6:::inh::D|
Imipenem|ok|Penicillin_binding_protein_4::STAAU:::D;PBPC::BACSU:inh::D;PBPA::ECOLI:inh::D;PBPB::ECOLI:inh::D;MRDA::ECOLI:inh::D|Beta_lactamase::KLEPN:sub::D;Q939N4,Q9L5C7,Q840M4:::sub::D;BLAT::ECOLX:sub::D;BLA1::ECOLX:sub::D;DPEP1:::sub::D||
Probucol|ok_inv|HEPS::::6.37:C;TAU::::5.15:C;EST1;ABCA1:::inh::D|||
Tiaprofenic_acid|ok|PGH1:::inh::D;PGH2:::inh::D|||
Lopinavir|ok|KCNH2::::5.07:C;Pol_polyprotein::9HIV1:inh::D|CP3A4,CP343,CP3A5,CP3A7:::inh:6.39,,,:DC;CP3A4:::inh:6.39:DC;CP2C8:::inh::D;CP2C9:::duo::D;CP2B6:::inh::D;CP2CJ:::inh::D;CP2D6:::inh::D|MDR1:::inh:5.77:DC;ABCBB:::sub::D;SO1B3:::inh::D;SO1B1:::inh::D|
Bacampicillin|ok_inv|PBPA::CLOPE:inh::D|||
Meticillin|ok_inv|PBPA::STRR6:inh::D;PBP3::STREE:inh::D;PBP2::STRR6:inh::D;PBP1B::STRR6:inh::D;PBP2A::STRR6:inh::D;MecA::STAAU:inh::D|||
Pivampicillin|ok|PBPA::CLOPE:inh::D|||
Pivmecillinam|ok|PBPA::CLOPE:inh::D|||
Tazobactam|ok|BLAT::ECOLX::7.77:C;AMPC::ENTCL::7.:C;BLA1::KLEPN::6.96:C;AMPC::MORMO::6.72:C;BLA1::ECOLX:inh:6.65:DC;AMPC::ECOLI::6.6:C;BLKPC::KLEPN::6.43:C;BLAC::STAAU::6.3:C;BLAC::BACLI::6.29:C;AMPC::PSEAE::6.09:C;AMPC::CITFR::6.03:C;BLO1::ECOLX::5.32:C;BLA1::ENTCL:inh::D;BLAT::SALTI:inh::D||S22A8:::inh::D;S22A6:::inh::D|
Ticarcillin|ok_inv_vet|PBP2A::STAAU:inh::D|||
Periciazine|ok_inv|LMNA::::8.2:C;CHLE::HORSE::6.64:C;ANDR::RAT::5.52:C;ACES::BOVIN::5.15:C;ANDR;ADA1B:::ant::D;ADA2A:::ant::D;DRD1:::ant::D|||
Deferasirox|ok_inv|Iron:::chel::D|CP1A2:::inh::D;CP2C8:::inh::D;UD19:::inh::D;UD13:::inh::D;UD11:::inh::D;CP3A4:::ind::D||
Valganciclovir|ok_inv|DNA:::cov::D||S15A1;S15A2;S6A14|
Hydroxychloroquine|ok|ACM2::::5.98:C;ADA1D::::5.63:C;TLR9:::ant::D;TLR7:::ant::D;DNA:::cov::D|CP2D6:::inh::D;CP3A4:::sub::D|SO1A2:::inh::D;MDR1:::inh::D|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Amyl_Nitrite|ok|ANPRA:::ago::D|ALDH2:::sub::D||
Erythrityl_tetranitrate|ok_exp_inv|ANPRA:::ago::D;ANPRB:::ago::D|||
Acepromazine|exp_vet|CP1A2::::5.8:C;CP2D6::::5.6:C;LEF::BACAN::5.6:C;PRIO::::5.3:C;LMNA::::5.25:C;TSHR::::5.1:C;ADA1B:::ant::D;ADA1A:::ant::D;5HT1A:::ant::D;5HT2A:::ant::D;DRD1:::ant::D;DRD2:::ant::D|||ALBU
Alverine|ok_inv|5HT1A:::ant::D|||
Molindone|ok|DRD2::RAT::7.48:C;5HT7R::::6.58:C;5HT2A::RAT::5.85:C;DRD1::RAT::5.8:C;ACM1;5HT2A:::ant::D;5HT1A:::ant::D;DRD2:::ant::D|||
Phenindamine|ok|HRH1::CAVPO::8.8:C;HRH1:::ant::D|||
Pheniramine|ok|HRH4:::ANT::D;NR1I3;HRH1:::ANT::D|||
Pipotiazine|ok_inv|DRD2:::ant::D;DRD1:::ant::D;5HT2A:::ant::D;5HT1A:::ant::D|CP3A4:::sub::D;CP2D6:::inh::D;CP2CJ:::sub::D|S22A1|ALBU
Thioproperazine|exp|ADA1B:::ant::D;ADA1A:::ant::D;5HT1A:::ant::D;5HT2A:::ant::D;DRD1:::ant::D;DRD2:::ant::D|||ALBU
Thiothixene|ok|5HT2A:::ant::D;DRD1:::ant::D;DRD2:::ant::D|CP2D6:::inh::D;CP1A2:::sub::D|S22A1|ALBU
Zuclopenthixol|ok_inv|DRD1:::ant::D;DRD5:::ant::D;DRD2:::ant::D;ADA1A:::ant::D;ADA2A:::ant::D;5HT2A:::ant::D;HRH1:::ant::D|CP2D6:::sub::D;CP3A4:::sub::D||
Isopropamide|ok_vet|LMNA::::5.45:C;CP2D6::::5.4:C;ACM4:::ant::D;ACM3:::ant::D|||
Pargyline|ok|AOFB:::inh:7.69:DC;TSHR::::6.9:C;CP3A4::::6.2:C;AOFB::RAT::5.55:C;AOFA:::inh:5.47:DC;ALDH2::RAT::5.25:C;AOFA::RAT::5.07:C;LMNA::::5.05:C|||
Lincomycin|ok_vet|RL10::SHIFL:inh::D|||
Etoricoxib|ok_inv|PGH2:::inh:7.09:DC;MK14::::6.28:C|CP2E1:::inh::D;CP2CJ:::inh::D;CP1A2:::sub::D;CP2D6:::inh::D;CP2C9:::inh::D;CP3A4:::inh::D||
5_O_phosphono_alpha_D_ribofuranosyl_diphosphate|ok_exp_inv|Hypoxanthine_guanine_phosphoribosyltransferase::TRYCR:::D;APT;Anthranilate_phosphoribosyltransferase::PECCA:::D;HPRT;PYRE::SALTY:::D;UCKL1|||
Sorbitol|ok|MASZ::ECOLI:::D;XYLA::ARTS7:::D;XYLA::ACTM4:::D;XYLA::STRRU:::D|||
Roflumilast|ok|PDE4D:::inh:9.57:DC;PDE4A:::inh:9.52:DC;PDE4B:::inh:9.4:DC;PDE4C:::inh::D|CP3A4:::sub::D||
Fumaric_Acid|exp_inv|TSHR::::5.4:C;FAAA;MAOM;FRDA::SHEON:::D;FRDA::SHEFR:::D;MDH::CHLAA:::D|||
Rutin|ok_exp_inv|ACES::::7.92:C;NMUR2::::5.92:C;LYAG::::5.5:C;MK01::::5.1:C;DPOLB::::5.05:C;ADA2A::::5.03:C;ADA2C::::5.02:C;CBR1;AK1C3|CP3A4:::inh::D||
Prasterone|ok_inv_nutra|SHBG::::7.84:C;GPBAR::::5.48:C;G6PD::::5.21:C;CBG::::5.:C;CHOD::BREST:::D;SDIS::PSEPU:::D;NR1I3:::act::D;NR1I2:::act::D;SGMR1:::ago::D;PPARA:::act::D;ST2B1;ST2A1;DHB1;ANDR:::ago::D;NMDA:::ago::D;GABAR:::ant::D;ESR2:::act::D;ESR1:::bin::D|CP3A7:::inh::D||
Cetrimonium|ok|MMAA2::MYCTU:::D;CMAS1::MYCTU:::D|||
Camphor|ok|AL1A1::::5.15:C;LMNA::::5.:C;TRPM8:::act::D;TRPA1:::inh::D;TRPV3:::ago::D;TRPV1:::ago::D;CPXA::PSEPU:::D|||
Dalfopristin|ok|VATD::ENTFC:inh::D|CP3A4:::inh::D||
Pantothenic_acid|ok_nutra_vet|COAA::ECOLI:::D|||
Propylene_glycol|ok_inv|B12_independent_glycerol_dehydratase::CLOBU:::D;FUCO::ECOLI:::D;CAS1::STRC2:::D;LINB::SPHJU:::D;F13A|||
D_glucose|ok_inv_vet||HXK1:::sub::D;HXK4:::sub::D|GTR1:::sub::D;GTR2:::sub::D;GTR3:::sub::D;GLUT4:::sub::D;GTR5:::sub::D;GTR6:::sub::D;GTR7:::sub::D;GTR8:::sub::D;GTR9:::sub::D;GTR10:::sub::D;GTR11:::sub::D;GTR12:::sub::D;SC5A1:::sub::D;SC5A2:::sub::D|
Taurine|ok_nutra|BLM::::7.9:C;GABR1:::ago::D;GABAR:::ago::D;GLRA3:::ago::D;GLRA2:::ago::D;NMDE2:::inh::D;GLRA1:::ago::D;CBH::CLOPE:::D;TAUD::ECOLI:::D|BAAT:::sub::D;TGM3L:::sub::D|S15A1:::sub::D;SC6A6:::sub::D;S36A1:::sub::D|
Cocarboxylase|ok_exp|MDLC::PSEPU:::D;POXB::LACPL:::D;DNA;ODP1::ECOLI:::D;PFOR::DESAF:::D;DCIP::ENTCL:::D;CEAS::STRCL:::D;TKT1::ECOLI:::D;ILVB::KLEPN:::D|||
Flufenamic_acid|ok|LMNA::::8.49:C;PGH2::::7.8:DC;AK1C3::::7.3:DC;TSHR::::6.7:C;AK1C2::::6.43:C;AK1BA::::6.12:C;AK1C1::::6.01:C;PERM::::5.74:C;PGH1::::5.65:DC;CP1A2::::5.4:C;HIF1A::::5.3:C;CP2C9::::5.:C;PPARG:::ago::D;PPARA:::act::D;ANDR||S22A6:::inh::D|TTHY::::5.54:DC
Calcipotriol|ok|VDR:::ant:9.51:DC|CP24A:::sub::D;PERM:::inh::D||
Isopropyl_alcohol|ok_inv|LMNA::::5.95:C;GUDD::ECOLI:::D;ENLYS::LAMBD:::D;POL::RSVSA:::D;MUTL::ECOLI:::D;DX39B;SAHH;PPA5;TNFA;Putative_deoxyribonuclease_YcfH::THEMA:::D;PRDX6;DCXR;Alr1529_protein::NOSS1:::D;CHIT1;Scaffolding_dockerin_binding_protein_A::CLOTM:::D;THER::GEOSE:::D;SAP3;PA2GA;MOP::DESGI:::D;GAG::SIVMK:::D;TRY2;Pectate_lyase::NIVIR:::D;RNAS1;KV401;SUBT::BACAM:::D;GDF5;GCH1;MTND;NUSG::AQUAE:::D;AZOR::ECOLI:::D;MCE1|||
Carbenoxolone|exp|DHI2::MOUSE::7.09:C;DHI1:::inh:7.08:DC;DHI1::MOUSE::6.97:C;HSD::STREX:::D|||
Aminobenzoic_acid|ok_exp|ACES::RAT::7.45:C;TSHR::::6.9:C;PHHY::PSEFL:::D;PHHY::PSEAE:::D|||
Tolrestat|out|ALDR::RAT::8.7:C;ALDR:::inh:8.:DC;AK1BA::::7.94:DC;ALDR::PIG::7.82:C;ALDR::BOVIN::7.48:C;AK1A1::PIG::6.27:C;AK1A1::::6.14:DC;AK1A1::RAT::5.92:C|||
Thymol|ok|LMNA::::6.1:C;TRPA1::::5.22:C|||
gamma_Aminobutyric_acid|ok_inv|BLM::::8.46:C;LMNA::::8.1:C;GBRP::RAT::7.89:C;GABR1::RAT::7.77:C;GBRA2::RAT::7.66:C;GBRA1::::7.6:C;GABR1::::7.6:DC;GBRG1::RAT::7.48:C;GBRR1::::6.57:C;GBRB2::::6.19:C;GBRG2::::5.82:C;SC6A1::RAT::5.79:C;GBRR2::::5.77:C;S6A11::RAT::5.7:C;GBRG2::RAT::5.64:C;GBRB3::::5.47:C;SC6A1::MOUSE::5.3:C;SC6A1::::5.3:C;S6A13::RAT::5.3:C;S6A11::::5.15:C;HDAC1::::5.09:C;S6A11::MOUSE::5.09:C;GBRA1::RAT::5.:C;GABR2;GATM||S36A1|
Vorinostat|ok_inv|HDAC6:::inh:9.:DC;HDAC1:::inh:8.89:DC;HDAC3:::inh:8.85:DC;HDAC2:::inh:8.8:DC;HDAC8::::8.26:DC;HDA11::::7.89:C;HDAC4::::7.8:C;HDAC9::::7.7:C;HDAC5::::7.48:C;HDAC7::::7.47:C;HDA10::::7.4:C;HDAC1::MOUSE::7.17:C;HDAC3::RAT::6.78:C;HDAH::ALCSD::6.52:C;NR0B1::::6.13:C;GLI1::MOUSE::5.65:C;NR1I2::RAT::5.6:C;PAX8::::5.34:C;Acetoin_utilization_protein::AQUAE:::D|||
Terlipressin|ok_inv|V1AR:::sti::D;V1BR;V2R:::ago::D|||
Fumagillin|exp|MAP2:::lig:9.2:DC|||
Cholic_Acid|ok|GPBAR::MOUSE::5.28:C;GPBAR::::5.22:DC;NR1H4;CBH::CLOPE:::D;Ferrochelatase;EST1;PA21B;CX7A1;CX6B1;CX6A2;COX8A;COX7C;COX7B;COX6C;COX5B;COX5A;COX3;COX2;COX1;COX41;FABP6;ERR3;ADH1G;HEMH||SO1B3:::sub::D;S22A7:::inh::D;S22A8:::inh::D;NTCP:::inh::D;MRP4:::inh::D;MRP3:::inh::D;SO1B1:::duo::D;MRP2:::ind::D;NTCP2:::duo::D;SO1A2:::duo::D;MRP1:::ind::D;MDR1:::ind::D;ABCBB:::duo::D|FABPL
Nicotinamide|ok_inv|SIR2::::5.92:C;FAAH1::RAT::5.48:C;TAU::::5.4:C;SIR3::::5.21:C;BST1;SIR5;PARP1:::bin::D;LDHA;TOXA::PSEAE:::D|CP3A4:::inh::D;CP2E1:::inh::D;CP2D6:::inh::D||
Fusidic_acid|ok_inv|ABCBB::RAT::5.66:C;MRP2::RAT::5.26:C;CAT3::ECOLX:inh::D;CAT::SALTI:inh::D;EFG::THETH:inh::D|UD11:::sub::D;CP3A4:::inh::D;CP2D6:::inh::D|SO1B1;ABCG2:::inh::D;MRP2:::inh::D;ABCBB:::inh::D|
Resveratrol|ok_exp_inv|LMNA::::8.3:C;NQO2::::7.27:DC;LUCI::PHOPY::7.23:C;AHR::RABIT::6.77:C;PK3CA::::6.6:C;PGH1::SHEEP::6.42:C;AOFA::::6.35:C;PK3CB::::6.3:C;PGH1:::inh:6.2:DC;TRPA1::RAT::6.12:C;PGH2:::inh:6.12:DC;ESR1::::6.11:DC;CAH9::::6.09:C;CAH14::::6.08:C;CAH12::::6.02:C;RORG::MOUSE::5.75:C;CAH1::::5.66:C;HD::::5.65:C;SC6A2::::5.64:C;NFKB2::::5.6:C;A4::::5.59:DC;CAH2::::5.56:C;CP2CJ::::5.52:C;PGH2::SHEEP::5.46:C;MTOR::::5.43:C;RAB9A::::5.4:C;ALR::::5.4:C;CAH13::::5.39:C;CAH7::::5.36:C;CAH4::::5.35:C;CAH5B::::5.33:C;CAH5A::::5.32:C;NF2L2::::5.27:C;NPC1::::5.25:C;TAU::::5.25:C;P53::::5.2:C;CP2C9::::5.15:C;CAH6::::5.09:C;SMN::::5.05:C;CAH3::::5.04:C;CAH15::MOUSE::5.03:C;PGDH::::5.:C;HIF1A::::5.:C;SYYC:::inh::D;FUBP2;AKT1:::inh::D;PPARG;PPARA;CBR1:::inh::D;GTR1;NR1I3;NR1I2;CLC14;MTR1B;MTR1A;SYUA;ITB3;ITA5;P4K2B;AHR;LOX5;LOX15;CSK21|CP3A4:::inh:6.22:DC;CP1A2:::inh:5.52:DC;CP1B1:::inh::D;CP1A1:::inh::D||ALBU;TTHY
Sucrose|ok_exp_inv|TS1R2;NTPPA::BACSU:::D;LYSC;NOSO::STAAW:::D;AMPC::ECOLI:::D;ACTS;ALGD::PSEAE:::D;SACB::BACSU:::D;SCRY::SALTM:::D;OCP::LIMMA:::D;RTCB;ATOX1;HMUO::CORDI:::D;Q939N4,Q9L5C7,Q840M4;Beta_lactamase::ECOLX:::D;AMYS::NEIPO:::D;Beta_glucosidase::STRSQ:::D|||
Pregnenolone|ok_exp|SHBG::::7.15:C;AMPC::ECOLI::6.5:C;CBG::::5.23:C;NR1I2;ST2B1|CP3A4:::sub::D|SOAT|
D_Methionine|ok_exp_inv|Transcriptional::VIBCH:::D;MAP2|||
Stanolone|ill_inv|ANDR::::10.3:DC;ANDR::RAT::9.57:C;ANDR::MOUSE::9.:C;SHBG::RAT::7.64:C;PRGR::RABIT::6.36:C;CBG::::5.92:C;MCR::RAT::5.68:C;GPBAR::::5.35:C;MCR;ESR1;DHB1|CP19A:::sub:6.66:DC;CP17A:::sub::D;CP11A:::sub::D|MDR1:::sub::D|SHBG::::9.74:DC
Piretanide|ok|LMNA::::8.4:C;HIF1A::::6.:C;UBP2::::5.1:C;AL1A1::::5.05:C;S12A1:::inh::D|||
Oxitriptan|ok_inv_nutra|5HT2C::::9.74:C;5HT1A::::9.04:C;5HT2B::::9.:C;5HT2A::::8.87:C;5HT7R::::8.67:C;5HT4R::RAT::8.01:C;LMNA::::7.4:C;5HT3A::RAT::6.8:C;NPSR1::::5.4:C;ACM1::RAT::5.35:C;TSHR::::5.3:C;AMPC::ECOLI::5.15:C;SYW2::DEIRA:::D|||
Lauric_acid|ok_exp|TSHR::::7.9:C;FFAR1::::6.12:C;PPARA;TLR4;LY96;PVDQ::PSEAE:::D;PA2GD;CO8G;TONB::ECOLI:::D;TRFL;FABF::ECOLI:::D;GLTP;VLDLR;PA2GA;HNF4A;POLG::HRV2:::D;POLG::HRV1A:::D;POLG::HRV16:::D;FABH::MYCTU:::D;SAP3;FHUA::ECOLI:::D;FABB::ECOLI:::D;ADHX|||ALBU
Glycolic_acid|ok_inv|GLYOX::BACSU:::D;G6PD|||
Pidolic_acid|ok_inv|LMNA::::8.25:C;AMY1;CSLB::PEDHD:::D;ANGI;AMY2B;CYCP::ALCXX:::D;CCL8;OREX;KRA52;Copper_containing_nitrite_reductase::ALCXX:::D;Endo::BACAG:::D;ADA28;CYC22::RHOPA:::D;TFF2;LV208;IGLC1;VEGFA|AMYP:::lig::DC||
Acetylcholine|ok_inv|ACM1::::8.96:DC;ACM5::::8.92:C;ACHB2::::8.77:C;ACM3::::8.49:DC;ACM2::::8.15:DC;ACHA4::RAT::8.12:C;ACM4::::8.:DC;ACHA2::RAT::7.96:C;ACM1::RAT::7.92:C;ACHA3::RAT::7.39:C;ACHA7::::6.3:DC;ACHA7::RAT::5.51:C;ACHP::LYMST::5.5:C;ACHD::TETCF::5.3:C;ACES||S22A1:::sub::D;S22A5:::inh::D|
Flavin_adenine_dinucleotide|ok|MEN1::::6.1:C;NDUA9:::cof::D;FRDA::SHEFR:::D;MRSD::BACSY:::D;FENR::ECOLI:::D;FENR::NOSS1:::D;AHPF::ECOLI:::D;DLDH::PSEFL:::D;DLDH1::PSEPU:::D;FkbI::STRHY:::D;Putative_acyl_CoA_dehydrogenase::THET2:::D;BENC::ACIAD:::D;PAMO::THEFY:::D;GSHR::PLAFK:::D;Dihydrolipoyl_dehydrogenase::NEIME:::D;AHPF::SALTY:::D;DH4C::PSEPU:::D;HDVD::CLOAM:::D;GLF::MYCTU:::D;LPDA::MYCTU:::D;CAMA::PSEPU:::D;Methylenetetrahydrofolate_reductase::THETH:::D;Phenol_2_hydroxylase_component_B::GEOTM:::D;HMP::ECOLI:::D;MURB::STAAW:::D;ALR;MURB::ECOLI:::D;ACOX1;ADRO;Oxidoreductase::BREST:::D;NB5R1;FRD2::SHEFN:::D;DLDH;CRYD::SYNY3:::D;NADB::ECOLI:::D;PHR::SYNP6:::D;PHR::ECOLI:::D;RNLS::PSESM:::D;DLDH::AZOVI:::D;Ferredoxin_reductase::PSES1:::D;AIFM1;ACDS::MEGEL:::D;ACAD8;FENR::AZOVI:::D;TRXR1;CYSJ::ECOLI:::D;DLD::ECOLI:::D;FENR::NOSSO:::D;DPYD;NAPE::ENTFA:::D;DMGO::ARTGO:::D;CHOD::BREST:::D;XDH;IVD;NQO2;TYTR::TRYCR:::D;MSOX::BACB0:::D;METF::ECOLI:::D;GSHR::ECOLI:::D;TRXB::ECOLI:::D;POXB::LACPL:::D;THYX::THEMA:::D;CHOD::STRS0:::D;NB5R3;FPRA::MYCTU:::D;GSHR;ERO1B;FRDA::SHEON:::D;PHHY::PSEFL:::D;NQO1;NOS1;PHHY::PSEAE:::D;XECC::XANP2:::D;FADH::ECOLI:::D;OXLA;ACADS;AOFA;PHR::THET8:::D;PUTA::ECOLI:::D;OXDA;ACADM;GCDH;NCPR;GLYOX::BACSU:::D;HMP::CUPNH:::D;GLF::ECOLI:::D|AOFB:::::DC||
Acetic_acid|ok|LCK::::6.19:C;FYN::::6.05:C||MOT1:::sub::D;SO2B1:::inh::D|
Propyl_alcohol|ok_exp|LYSC|||
Stearic_acid|ok_exp|PPARA::::5.96:DC;PPARD::::5.22:C;TSHR::::5.:C;PA2GD|||ALBU;FABPH
Oteracil|ok|LMNA::::6.55:C|||
Flavin_mononucleotide|ok_inv|IDI2::THET2:::D;FPRA::MOOTA:::D;NFSB::ENTCL:::D;SGK1;FLAV::HELPJ:::D;AZR::BACSU:::D;MDLB::PSEPU:::D;PADL::ECO57:::D;NRDI::BACSU:::D;tRNA_dihydrouridine_synthase::THEMA:::D;MOXC::BACSU:::D;Uncharacterized_protein::STRMU:::D;FLAV::SYNE7:::D;FLAV::DESVH:::D;FLAV::NOSS1:::D;AROC::HELPY:::D;AZOR::ECOLI:::D;EPID::STAEP:::D;AZOR::SALTY:::D;Pentaerythritol_tetranitrate_reductase::ENTCL:::D;PYRD;DPYD;PYRD::ECOLI:::D;NOS1;NFSA::ECOLI:::D;RIFK;FRA1::ALIFS:::D;PNPO;HAOX1;BLVRB;PYRDA::LACLC:::D;FADH::ECOLI:::D;AROC::STRR6:::D;NFSB::ECOLI:::D;FLAV::CLOBE:::D;PDXH::ECOLI:::D;GLTS::SYNY3:::D;Phenazine_biosynthesis_protein::PSEAI:::D;COAC;Nitroreductase_family_protein::BACCR:::D;FMNB::DESVM:::D;NOX::THET8:::D;IDI2::BACSU:::D;FLAV::ECOLI:::D;NQOR::DEIRA:::D;HAOX2;PHZG::PSEFL:::D;KS6A4;FRP::VIBHA:::D;Morphinone_reductase::PSEPU:::D;Riboflavin_biosynthesis_protein::THEMA:::D;ROO::DESGG:::D;DHTM::METME:::D|NCPR:::lig::DC||
Phenol|ok_exp|CAH3::::5.57:C;CAH2::::5.26:C;CAH9::::5.06:C;CAH12::::5.04:C;CAH4::::5.02:C;CAH1::::5.:C;AGAL::::5.:C;ALBU;COBT::SALTY:::D;ENLYS::BPT4:::D;THER::GEOSE:::D|||
Glutathione_disulfide|ok_exp_inv|GSHR;GSTM2|||
Brivudine|ok_inv|KITH::::7.:C;KITH::HHV1::6.62:C;KITH::HHV1S::6.52:C;CYSP::TRYCR::5.5:C;KITH::HHV11:::D|||
Hemin|ok_inv||||
Oxyphenbutazone|ok_out|RORG::MOUSE::5.35:C;PA2GE||S22A6:::inh::D|ALBU
Tiratricol|inv|THB::::10.39:DC;THA::::9.85:C;THB::RAT::9.82:C;SO1C1::MOUSE::5.67:C;CP2C9::::5.3:C;HIF1A::::5.2:C;HCD2::::5.:C|||
Methylcobalamin|ok_exp_inv|METH::ECOLI:::D|||
Ribostamycin|ok_exp|RS12::ECOLI:::D;PDIA1;AAC6::SALEN:::D|AAC2::MYCTU:sub::DC||
Deoxycholic_acid|ok|GPBAR::::5.9:DC;GSTP1;NR1H4;COX2::RHOSH:::D;COX1::RHOSH:::D;ACRB::ECOLI:::D;ALDA::ECOLI:::D;CBH::CLOPE:::D;EFL1;Cytochrome_C::GEOSN:::D;SDIS::PSEPU:::D||NTCP2:::inh:5.2:DC;NTCP:::sub::D;SO1A2:::inh::D;ABCBB:::ind::D|
Tromethamine|ok|LMNA::::6.45:C;PGS2;6PGL::THEMA:::D;VEGFA;BIOB::ECOLI:::D;DCAM;CHTB::VIBCH:::D;NEIL1;Y1317::HAEIN:::D;DPS::AGRFC:::D;NLPI::ECOLI:::D;CANT1;CYC4::PSEST:::D;ALYS::STRPN:::D|||
Doconexent|ok_inv|OXER1::::5.7:C;PGH2::SHEEP::5.01:C;SRBP1:::inh::D;RXRG:::act::D;RXRB:::act::D;RXRA:::act::D;PPARG:::lig::D;PPARA:::lig::D|CP2C9:::inh::D||FABP7
Propanoic_acid|ok_vet|ALR::GEOSE:::D;2::PSEFL:::D;GEPH;PRXC::PSEFL:::D|||FABP4
Phenacetin|out|MEN1::::5.:C;PGH1|CP1A2:::sub:5.:DC;CP3A4:::sub::D;CP2E1:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP2A6:::sub::D;CP2AD:::sub::D;CP1A1:::sub::D;CP2D6:::sub::D|S22A6:::inh::D|
Benzoic_acid|ok_inv|LEF::BACAN::5.9:C;OXDA::::5.7:DC;TSHR::::5.:C;S15A1;COCE::RHOSM:::D;ELBP::ECOLX:::D;PRDX5;Replication_protein::PSESX:::D;CHQB::NOCSI:::D;NFSB::ENTCL:::D;PRXC::KITAU:::D;2::PSEFL:::D;RAB9A;CLCA::RHOOP:::D;RIDA;PPTA::ECOLI:::D;MALT::ECOLI:::D;OXYR::ECOLI:::D||MOT1;S22A8:::inh::D;SO2B1:::inh::D|
Palmitic_Acid|ok|PPARA::::5.82:DC;TLR2::::5.3:C;PPARD::::5.13:C;LALBA;MYP2;PPT1;S14L2;OPSD;Y1468::THEMA:::D;TPPC3;CP2C8;Lipid_binding_protein::GEOSE:::D;HNF4G;PAEP|||FABP4::::6.47:DC;FABP5::::6.1:DC;FABPI::::5.77:DC;FABPH::::5.59:DC;ALBU
Hexamidine|exp|THRB::::6.65:C;ST14::::6.03:C;QACR::STAAU:::D;QACR::STAHA:::D|||
Formaldehyde|ok_vet|DAC::STRSR:::D|||
Eucalyptol|exp_nutra||||
Urea|ok_inv|LMNA::::6.1:C;DYR::ECOLI:::D;MSRP::ECO57:::D;CTNB1;POLS::EEVVT:::D;CAH2;ARGI1||UT1:::sub::D;UT2:::sub::D|
D_Serine|ok_exp|BLM::::8.6:C;NMDZ1::RAT::6.8:C;DECO::BPP21:::D;SPB3;NMDZ1;GLRA1||S6A14;MOT10:::inh::D|
Ergosterol|ok_exp||||
Fotemustine|inv|TRXR1|||
Berberine|ok_inv|ACES::::7.:C;ACES::ELEEL::6.43:C;CHLE::::5.96:C;HIF1A::::5.6:C;CP2D6::::5.6:C;CP1A2::::5.3:C;BIRC5;QACR::STAHA:::D|||
Nicotinyl_alcohol|exp||||
Pyrophosphoric_acid|ok_exp|IDI::ECOLI:::D;ISPA::ECOLI:::D;FHUA::ECOLI:::D;KTHY::MYCTU:::D;NADE::ECOLI:::D;PURA::SHIFL:::D|||
Valpromide|exp|LIMA::RHOER:::D|||
Fructose|ok_exp|LAMB::ECOLI:::D;FHIT|||
Dequalinium|ok_inv|LMNA::::6.1:C;CP3A4::::5.8:C;ACM1::RAT::5.75:C;HIF1A::::5.7:C;RORG::MOUSE::5.65:C;TAU::::5.5:C;FFP::BACIU::5.35:C;TPO::::5.3:C;MTOR::::5.13:C;TSHR::::5.1:C;HD::::5.1:C;CP1A2::::5.:C;CP2D6::::5.:C;KCMA1:::inh::D;CNGA1:::inh::D;XIAP:::ant::D;QACR::STAHA:::D;ACRB::ECOLI:::D|||
Didecyldimethylammonium|ok_exp|CMAS2::MYCTU:::D|||
Oleic_Acid|ok_inv_vet|PPARG:::lig::D;RXRA;PPARD;PPARA;MYP2;FABP::SCHMA:::D;GLTP|||VTDB;ALBU;FABPL;FABPH;FABP4;FABP7
Citric_acid|ok_nutra_vet|AROQ::HELPY::5.6:C;AROQ::STRCO::5.14:C;BLAC::BACLI:::D;ECP;GNMT;IDH::BACSU:::D;RNAS1;PDC::ZYMMO:::D;SRC;PCAB::PSEPU:::D;PDE5A;Glycerol_uptake_operon_antiterminator_regulatory_protein::THEMA:::D;HS3SA;ENLYS::BPP1:::D;CISY;ITPA;ALDR;GUAA::ECOLI:::D;SYW::GEOSE:::D;RPIA::HAEIN:::D;BHMT1;POLOX::ECOLI:::D;TN13B;UCK2;Glyoxalase_family_protein::BACCR:::D;BLA2::BACCE:::D;Glucose_1_phosphate_thymidylyltransferase::PSEAE:::D;ANGI;APT;FTSZ::MYCTU:::D;PGFS::TRYBB:::D;PRPC::ABDS2:::D;GLN1B,GLN1B::MYCTO,MYCTU:::D;RIR2::MYCLE:::D;CO8G;NUSB::THEMA:::D;NADD::SHIFL:::D;Signal_recognition_particle_receptor_FtsY::THEMA:::D;FBPA::SERMA:::D;PKHA1;LSM6;RTCA::ECOLI:::D;Citrate_synthase::THETH:::D;Putative_stringent_starvation_protein_A::YERPE:::D;BFRA::THEMA:::D;Riboflavin_biosynthesis_protein::THEMA:::D;CAPSH::ADE02:::D;CBPB1;RL4::THEMA:::D;N5_carboxyaminoimidazole_ribonucleotide_mutase::ACEAC:::D;MDHM;FIB12::BPT4:::D;TEV1::BPT4:::D;INVA::YERPS:::D;HGS;Cytochrome_c_peroxidase::MARHY:::D;NANH::MICVI:::D;TRPA::THET2:::D;DXR::ECOLI:::D;CTDS1;MIF;OXLA;POL::RSVSA:::D;NFSB::ECOLI:::D;6PGL::THEMA:::D;FUMC::ECOLI:::D;MOBA::ECOLI:::D;ALKH::ECOLI:::D||SO2B1:::inh::D|
Inosine|exp_inv|DEOD::ECOLI:::D;PNPH;IAG_nucleoside_hydrolase::TRYVI:::D|XDH:::sub_ind::D|S28A3|
Carbocisteine|ok_inv|GSTP1|||
Taurocholic_acid|ok_exp|GPBAR::::5.31:C;NTCP::RAT::5.22:C;NR1H4;FABP6;CEL||NTCP:::sub:5.28:DC;XCT;SO1B3:::sub::D;OSTB:::sub::D;OSTA:::sub::D;MOT1:::sub::D;SO2B1:::sub::D;ABCG2:::inh::D;SO3A1:::inh::D;SO1C1:::inh::D;ABCCB:::inh::D;SO4A1:::inh::D;S22A8:::inh::D;MRP7:::inh::D;S22A6:::inh::D;MDR1:::inh::D;MRP4:::inh::D;MRP3:::inh::D;SO1B1:::duo::D;MRP2:::ind::D;NTCP2:::sub_ind::D;SO1A2:::duo::D;MRP1:::duo::D;ABCBB:::sub_ind::D|
Meglutol|exp|HMDH::::7.63:DC|||
Lactic_acid|ok_vet|P53::::7.6:C;NimA_related_protein::DEIRA:::D;PUTA::ECOLI:::D||MOT4:::sub::D;SO2A1:::inh::D;MOT10:::inh::D;MOT1:::inh::D;SO2B1:::inh::D;MOT2:::inh::D|
Mercuric_iodide|exp|ST2A1|||
Lactose|ok_exp_inv|GL6D1;GLTP;ETXB::STAAU:::D;NANH::MICVI:::D;Beta_xylanase::STROI:::D;XYNA::STRLI:::D;BGAL::ECOLI:::D;TETX::CLOTE:::D;LEG3|||
Cholesterol|ok_inv|LMNA::::5.2:C;CLC4E:::lig::D;VDR;NR1I3;RORA||MDR1:::inh:5.09:DC;ABCG2:::ind::D|
Niflumic_acid|exp|KPYM::::7.6:C;TTHY::::6.59:C;PGH2:::inh:6.04:DC;PGH1::::5.97:DC;GPR35::::5.95:C;NFKB1::::5.65:C;CP1A2::::5.3:C;HIF1A::::5.2:C;CP3A4::::5.1:C;PA24A;CLCKA:::ind::D;PA21B:::inh::D|UD19:::inh::DC|MOT1:::inh::D;MOT2:::inh::D|
Gluconolactone|ok_exp|LMNA::::6.1:C;LPH|||
Latamoxef|ok_inv|DACB::ECOLI:inh::D;PBPB::ECOLI:inh::D;PBPA::ECOLI:inh::D;PBPC::BACSU:inh::D|||
Trioxsalen|ok|KDM4E::::6.55:C;AA2AR::::6.13:C;AOFA::::6.08:C;CP1A2::::6.:C;5HT2C::::5.91:C;AL1A1::::5.45:C;CP3A4::::5.4:C;MK01::::5.2:C;DNA:::cov::D|||
Thiotepa|ok_inv|HBB::::5.6:C;PGDH::::5.:C;LMNA::::5.:C;DNA:::cov::D|CP2B6:::inh:5.66:DC;CHLE:::inh::D;CP3A4:::sub::D||
Estriol|ok_inv_vet|ESR2:::ago:9.9:DC;ESR1:::ago:9.32:DC;SHBG::::6.63:DC;SC6A4::::5.26:C;LOX15::RABIT::5.06:C;SO1A1::RAT::5.01:C;CBG::::5.:C||MDR1:::sub_ind::D;SO1A2:::inh::D|
Estrone_sulfate|ok|SO1B1::::7.34:C;MRP1::::6.35:C;SO1A1::RAT::5.89:C;STS::::5.12:C;S22A8::RAT::5.04:C;ESR2:::ago::D;ESR1:::ago::D|CP2C9:::inh::D;CP1A2:::sub::D;CP3A4:::sub::D|S47A2:::sub::D;S47A1:::sub::D|ALBU;SHBG
Quinestrol|ok|LMNA::::6.95:C;STRP::STRP1::5.58:C;ESR1:::ago::D|||
Fleroxacin|exp|KDM4E::::5.5:C;PARC::HAEIN:inh::D;GYRA::HAEIN:inh::D;TOP2A:::inh::D|||
Aniracetam|exp|BLM::::8.4:C;RECQ1::::6.65:C;TAU::::6.25:C;THB::::5.95:C;CP2CJ::::5.7:C;CP2C9::::5.2:C;GRIA3;GRIA2;DRD2;5HT2A|||
Aldosterone|exp_inv|MCR::::9.74:DC;MCR::RAT::7.37:C;CBG::::6.28:C;SHBG::::5.32:C;GCR|CP3A4:::sub::D;CP17A:::ind::D;C11B2:::sub::D;C11B1:::sub::D|SO1A2:::inh::D;S22A5:::inh::D;MDR1:::sub_ind::D|
Carboxin|ok_exp|MK01::::5.5:C;HCD2::::5.4:C;SDHA|||
Choline_alfoscerate|exp_inv|AMPC::ECOLI::6.25:C;SAP3|||
Hesperidin|ok_inv|CAC1B::::5.02:C;AURKB|||
Iodipamide|ok|TSHR::::5.2:C|||ALBU:::bin::D
Nimesulide|ok_out|PGH2:::inh:9.:DC;PTGES::MOUSE::8.15:C;PGH2::MOUSE::8.15:C;CP2D6::::7.3:C;CP2CJ::::7.1:C;TSHR::::7.:C;LMNA::::6.9:C;PGH2::SHEEP::6.4:C;CP19A::::6.17:C;PGH1::::5.91:C;PGH1::MOUSE::5.78:C;PERM::::5.68:C;HIF1A::::5.5:C;CP2C9::::5.5:C;CP1A2::::5.4:C;AGAL::::5.4:C;PGH1::SHEEP::5.21:C;PTGES::::5.:C;TRFL;PA2GE|CP3A4:::sub::D||
Suramin|inv|P2Y11::::6.95:C;SIR1::::6.52:C;P2RX1::RAT::6.:C;SIR2::::5.96:C;NR1I2::::5.89:C;PRKDC::::5.77:C;SIR5:::inh:5.7:DC;RECQ1::::5.6:C;PFKA::TRYBB::5.52:C;P2RX3::::5.52:C;UBP2::::5.48:C;P2RX2::RAT::5.4:C;P2Y12::RAT::5.4:C;P2RX5::RAT::5.4:C;TYDP1::::5.35:C;ANM1::::5.27:C;HCD2::::5.1:C;VCP::VACCW:::D;PA2GA:::inh::D;THRB:::inh::D;RYR1:::ago::D;FSHR:::ant::D;P2RY2:::ant::D|PA24A:::inh::D;ARSA:::inh::D||
Bifonazole|ok_inv|CP17A::::7.25:C;CP51A::::6.47:C;HS90A::::5.97:C;HIF1A::::5.9:C;RORG::MOUSE::5.5:C;MEN1::::5.5:C;ATG4B::::5.07:C;PA21B::::5.05:C;AL1A1::::5.05:C;CP2B6;CP51::CANAL:inh::D|CP3A4:::inh:7.:DC;CP2E1:::inh::D;CP19A:::inh::D||
Benoxaprofen|ok_out||||
Bithionol|ok_out|MK14::::6.5:C;MK01::::6.41:C;AA3R::::6.33:C;ADA2B::::6.25:C;EGFR::::6.21:C;ADA2C::::6.2:C;AA2AR::::6.18:C;LOX12::::6.15:C;NR1I2::::6.:C;SC6A2::::5.91:C;ADA2A::::5.84:C;DRD3::::5.84:C;NK2R::::5.81:C;SC6A3::::5.76:C;THAS::::5.74:C;S22A2::::5.72:C;MCL1::::5.72:C;ERBB2::::5.67:C;OPRM::::5.65:C;LCK::::5.65:C;LEF::BACAN::5.5:C;LMNA::::5.5:C;5HT1A::RAT::5.5:C;S22A1::::5.41:C;ESR1::::5.4:C;5HT2B::::5.36:C;5HT2C::::5.34:C;HIF1A::::5.3:C;S47A1::::5.28:C;S22A3::::5.26:C;S47A2::::5.18:C;ESR2::::5.09:C;TAU::::5.:C;HD::::5.:C|||
Clioquinol|ok_vet_out|CP1A2::::7.5:C;HIF1A::::7.4:C;LMNA::::7.:C;RORG::MOUSE::6.45:C;LOX12::::6.15:C;HS90A::::5.94:C;CAH15::MOUSE::5.63:C;COMT::RAT::5.32:C;P53::::5.3:C;OPRK::::5.24:C;HD::::5.:C|||
Dantron|ok_out|TSHR::::5.7:C;MK01::::5.5:C;TAU::::5.3:C;LMNA::::5.:C;RORG::MOUSE::5.:C|||ALBU
Metamizole|ok_out|PGH1|CP3A4:::ind::D;CP2B6:::ind::D||
Iproniazid|out|AOFA::RAT::5.3:C;AOFB::RAT::5.12:C|AOFB:::inh:5.71:DC;AOFA:::inh:5.59:DC;CP2C9:::inh::D;CP2D6:::inh::D||
Methapyrilene|out||||
Nialamide|ok_out|CYSP::TRYCR::6.7:C;END4::ECOLI::5.25:C;TSHR::::5.2:C;LMNA::::5.15:C;CP2D6::::5.1:C;KDM4E::::5.05:C;CP2CJ::::5.:C;CP2C9::::5.:C;COMT;AOFA;AOFB|||
Nomifensine|ok_out|SC6A2::::8.3:DC;SC6A3::::8.:DC;SC6A3::RAT::7.59:C;DRD5::RAT::7.32:C;SC6A4::RAT::6.08:C;SC6A4::::5.85:DC;VMAT2;PERM;AOFA;AOFB|||A1AG1
Oxeladin|ok_out||||
Oxyphenisatin|inv_out||||
Phenolphthalein|ok_out|LMNA::::7.6:C;TYSY::::5.92:C;TYSY::ENTFA::5.85:C;LEF::BACAN::5.6:C;CP3A4::::5.4:C;TYSY::LACCA::5.33:C;TYSY::ECOLI::5.33:C;GPR55::::5.18:C;SHBG;ESR1:::ago::D;NR1I3;NR1I2;UD19|||
Prenylamine|ok_out|KCNH2::::7.19:C;CAC1C::RAT::6.68:C;SCN1A::::6.52:C;CALM::BOVIN::6.3:C;CAC1C::CAVPO::5.91:C;SCN5A::::5.6:C;MYLK2:::inh::D;CALM1|CP3A4:::sub::D||
Thenalidine|ok_out||||
Urethane|ok_out||AOXA:::sub::D;PERM:::ind::D;PA24A:::sub::D||
Zomepirac|out|PD2R2|CP3A4:::sub::D||ALBU
Buformin|inv_out|LMNA::::5.5:C||S22A1:::sub::D|
Tienilic_acid|out|ALDR::RAT::5.49:C|CP2C9:::inh:5.37:DC||
Zimelidine|ok_out|SC6A4::RAT::5.35:C;AOFA:::inh::D;AOFB:::inh::D;SC6A4|CP3A4:::inh::D|MDR1:::inh::D|
Methaqualone|ill_out|LMNA::::6.5:C|CP3A4:::sub::D||
Rapacuronium|ok_out|ACM2:::ant::D|||
Maraviroc|ok_inv|CCR5:::ant:9.7:DC;CCR5::MACMU::9.62:C|CP3A4:::sub::D||
Amineptine|ill_out|SC6A2;SC6A4|||
Clofedanol|ok_out|HRH1:::ant::D|||
Cyclandelate|ok|EST1;CA2D1:::inh::D|CP3A4:::sub::D||
Cyproterone_acetate|ok_inv|AA1R::RAT::9.12:C;ANDR:::ant:7.85:DC;ANDR::RAT::7.51:C;GCR::::6.99:C;AA2BR::RAT::6.47:C;OPRM::::6.05:C;RORG::MOUSE::5.85:C;KLK3|CP3A4:::inh:5.6:DC;CP19A:::inh::D||
Debrisoquine|ok_inv|SC6A2:::ind::D|CP1A1:::sub::D;CP2D6:::sub::D|MDR1:::sub::D|
Flunarizine|ok|LMNA::::8.49:C;SGMR1::::8.:C;HRH1:::ant:7.74:DC;ADA2C::::7.49:C;DRD3::::7.48:C;SCN2A::RAT::7.28:C;CA2D1::RAT::7.1:C;CP2J2::::7.:C;5HT2A::::6.94:C;DRD2::::6.93:C;ADA2A::::6.66:C;DRD2::RAT::6.64:C;SC6A4::::6.58:C;ACM3::::6.5:C;5HT2C::::6.45:C;ADA1A::RAT::6.36:C;SC6A3::::6.33:C;KCNH2::::6.3:C;CAC1G:::inh:6.28:DC;ADA1D::::6.27:C;SCN1A::::6.22:C;ADA1B::RAT::6.22:C;5HT2B::::6.16:C;ACM1::::6.15:C;ACM4::::6.1:C;ACM5::::6.1:C;CAC1I:::inh:6.08:DC;ADA2B::::6.06:C;SC6A2::::5.88:C;CAC1B::::5.78:C;DRD1::::5.71:C;OPRM::::5.67:C;CNR1::::5.62:C;5HT1A::RAT::5.61:C;AA3R::::5.53:C;CAC1H:::inh:5.44:DC;CALM1|CP2D6:::sub:5.1:DC;CP3A4:::sub::D;CP2A6:::sub::D;CP1A2:::sub::D;CP1A1:::sub::D;CP2C9:::sub::D||
Fluspirilene|ok_inv|5HT2B::::6.82:C;OPRX::::6.3:C;LMNA::::6.:C;5HT6R::::5.93:C;GLRA1::::5.92:C;CP2D6::::5.8:C;KCNH2::::5.64:C;LYAG::::5.3:C;MEN1::::5.2:C;CP2CJ::::5.1:C;NPSR1::::5.1:C;DNAB::MYCTU::5.01:C;XBP1::::5.:C;TAU::::5.:C;NFKB1::::5.:C;CCG1:::inh::D;5HT2A:::ant::D;DRD2:::ant::D|CP3A4:::sub:5.2:DC||
Mepenzolate|ok|ACM1:::ant::D;ACM3:::ant::D|||
Tetrabenazine|ok_inv|VMAT2::BOVIN::8.4:C;VMAT2::RAT::8.12:C;DPOLB::::5.4:C;DRD2:::inh::D;VMAT2:::inh::D|CBR1:::sub::D;CP2D6:::sub::D||
Ixabepilone|ok_inv|TBB3:::inh::D|CP3A4:::inh::D||
Celiprolol|ok_inv|5HT1A::RAT::5.05:C;ADA2C:::ant::D;ADA2B:::ant::D;ADA2A:::ant::D;ADRB3:::ago::D;ADRB2:::ago::D;ADRB1:::ant::D|CP2D6:::sub::D||
Roxadustat|inv|EGLN1::::6.23:DC;FTO::::5.01:C;EGLN3;EGLN2|||
Cediranib|inv|KIT:V559D:::9.57:C;KIT:V559D-V654A:::9.51:C;KIT:V559D-T670I:::9.49:C;PGFRB::::9.49:C;KIT::::9.42:C;PGFRA::::9.39:C;KIT:L576P:::9.27:C;VGFR1::::9.13:C;VGFR2::::9.:DC;DDR1::::8.77:C;VGFR3::::8.52:C;STK35::::8.27:C;RET::::8.21:C;RET:M918T:::8.12:C;FGFR3::::7.9:C;CSF1R::::7.89:C;SLK::::7.8:C;ABL1:T315I:::7.7:C;STK10::::7.64:C;FGFR1::::7.6:C;FGFR2::::7.46:C;FGFR3:G697C:::7.46:C;EPHA6::::7.44:C;ABL1:H396P:::7.41:C;PTK6::::7.4:C;DDR2::::7.32:C;SRC::::7.3:C;M4K5::::7.3:C;ABL1:Y253F:::7.26:C;ABL1:M351T:::7.25:C;LYN::::7.2:C;ABL1:E255K:::7.19:C;LCK::::7.17:C;ABL1:Q252H:::7.11:C;ABL1::::7.11:C;FRK::::7.1:C;EGFR:G719S:::7.08:C;KIT:A829P:::7.01:C;RIPK2::::7.01:C;EGFR:L861Q:::6.92:C;BLK::::6.92:C;EGFR:L858R:::6.85:C;TIE2::::6.85:C;EGFR:G719C:::6.82:C;ERBB3::::6.74:C;EPHB6::::6.66:C;EGFR::::6.64:C;M3K19::::6.6:C;YES::::6.59:C;ABL1:F317L:::6.55:C;TIE1::::6.54:C;UFO::::6.5:C;MET::::6.43:C;KIT:D816V:::6.41:C;ERBB2::::6.4:C;FYN::::6.3:C;ERN1::::6.29:C;STK33::::6.27:C;MINK1::::6.27:C;M4K2::::6.27:C;MET:Y1235D:::6.25:C;MET:M1250T:::6.24:C;HCK::::6.23:C;EPHA7::::6.21:C;ABL2::::6.14:C;TNIK::::6.09:C;KIT:D816H:::6.09:C;TYRO3::::6.08:C;FGFR4::::6.07:C;M4K1::::6.04:C;RON::::6.:C;LTK::::6.:C;FER::::6.:C;FGR::::5.96:C;EPHB4::::5.96:C;ERBB4::::5.9:C;M4K4::::5.9:C;AURKB::::5.9:C;KSYK::::5.9:C;ABL1:F317I:::5.89:C;EGFR:T790M:::5.89:C;MP2K5::::5.82:C;ACV1B::::5.82:C;TAOK1::::5.8:C;GAK::::5.77:C;TGFR1::::5.77:C;ACVR1::::5.7:C;KPCD2::::5.7:C;PLK4::::5.7:C;M4K3::::5.7:C;SIK2::::5.68:C;AURKC::::5.68:C;FLT3:K663Q:::5.64:C;ALK::::5.64:C;CHK2::::5.6:C;MERTK::::5.59:C;KC1E::::5.55:C;E2AK1::::5.51:C;MP2K2::::5.51:C;EPHA3::::5.43:C;RET:V804M:::5.42:C;STK3::::5.4:C;STK4::::5.37:C;BTK::::5.37:C;STK26::::5.35:C;TAOK3::::5.3:C;KCC2B::::5.3:C;EPHA1::::5.28:C;EPHA8::::5.28:C;TAOK2::::5.23:C;EGFR:L858R-T790M:::5.13:C|||
Febuxostat|ok|XDH::BOVIN::9.92:C;XDH:::inh:8.9:DC;XDH::RAT::8.4:C|||
Dronedarone|ok|KCNH2:::inh:6.5:DC;CAC1C::CAVPO::6.4:C;THA:::inh::D;KCND3:::inh::D;NAC1:::inh::D;KCJ12,KCJ14,KCNJ2,KCNJ4:::inh::D;KCNQ1:::inh::D;KCNJ3:::inh::D;SCN5A:::inh::D;KCNK2:::inh::D;CACB4:::inh::D;CACB3:::inh::D;CACB2:::inh::D;CACB1:::inh::D;CAC1S:::inh::D;CAC1F:::inh::D;CAC1D:::inh::D;CAC1C:::inh::D;ADRB1:::ant::D;ADA2C:::ant::D;ADA2B:::ant::D;ADA2A:::ant::D;ADA1D:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D|CP2J2:::inh::D;CP3A5:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D|S22A8:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;S22A1:::inh::D;S22A2:::inh::D;MDR1:::inh::D|ALBU:::bin::D
Nebivolol|ok_inv|KCNH2::::6.5:C;SCN5A::::5.2:C;ADRB3:::ago::D;ADRB2:::ant::D;ADRB1:::ant::D|CP2CJ:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D||ALBU:::bin::D
Huperzine_A|ok_exp|ACES::RAT::7.09:C;ACES:::inh:6.22:DC|||
Omacetaxine_mepesuccinate|ok_inv|RL3:::ant::D;RL2::HALMA:ant::D|||
Nilotinib|ok_inv|ABL1:::inh:9.48:DC;DDR1::::8.96:C;DDR2::::8.7:C;CAH2::::8.39:C;ABL1:H396P::inh:8.31:DC;ABL1:Q252H::inh:8.:DC;M3K20::::7.96:C;ABL1:F317L::inh:7.92:DC;ABL1:Y253F::inh:7.89:DC;ABL1:M351T::inh:7.89:DC;KIT:::ant:7.83:DC;PGFRB::::7.8:C;ABL1:F317I::inh:7.74:DC;KIT:L576P::ant:7.66:DC;ABL2::::7.59:C;ABL1:E255K::inh:7.56:DC;CAH1::::7.53:C;MK11::::7.44:C;EPHA8::::7.43:C;CAH9::::7.38:C;CSF1R::::7.35:C;KIT:A829P::ant:7.34:DC;KIT:V559D::ant:7.34:DC;LCK::::7.33:C;PGFRA::::7.15:C;CAH15::MOUSE::7.1:C;FRK::::7.07:C;LYN::::7.:C;CAH7::::7.:C;EPHA3::::6.96:C;KCNH2::::6.9:C;KIT:V559D-T670I::ant:6.82:DC;MP2K5::::6.72:C;ABL1:G250E::inh:6.67:DC;CAH14::::6.65:C;EPHA2::::6.64:C;KIT:V559D-V654A::ant:6.59:DC;CAH12::::6.52:C;FGR::::6.49:C;EPHA4::::6.48:C;TNI3K::::6.44:C;NQO2::::6.42:C;HCK::::6.41:C;MK08::::6.35:C;CAH3::::6.35:C;CAH4::::6.35:C;MK14::::6.34:C;CAH6::::6.34:C;NTRK2::::6.31:C;BLK::::6.3:C;EPHB6::::6.3:C;KIT:D816H::ant:6.27:DC;BRAF:V600E:::6.24:C;EPHA1::::6.23:C;NTRK3::::6.22:C;EPHB2::::6.19:C;EPHA6::::6.19:C;ABL1:T315I::inh:6.18:DC;EPHB4::::6.14:C;KIT:D816V::ant:6.11:DC;CDPK1::PLAF7::6.1:C;RET::::6.06:C;M4K1::::6.05:C;MRCKB::::6.04:C;TIE1::::6.:C;TIE2::::6.:C;EPHB3::::6.:C;YES::::5.96:C;RET:M918T:::5.96:C;RAF1::::5.96:C;EPHB1::::5.89:C;FYN::::5.8:C;TAOK3::::5.77:C;BRAF::::5.77:C;SRC::::5.72:C;EPHA5::::5.72:C;MK10::::5.7:C;CLK1::::5.68:C;CSK::::5.62:C;TAOK1::::5.33:C;CAC1C::::5.33:C;CAH13::MOUSE::5.33:C;CAH5A::::5.26:C;MK09::::5.24:C;STK10::::5.17:C;CLK4::::5.15:C;PI42C::::5.06:C;FLT3::::5.02:C|CP2B6:::ind::D;CP2D6:::inh::D;CP2C9:::inh::D;CP2C8:::duo::D;CP3A4:::inh::D|SO1B1:::inh::D;UD11:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|
Lorcaserin|ok|5HT2B::::8.89:C;5HT2A::::8.89:C;5HT2C::::8.74:DC;5HT2C::CANLF::7.79:C;SC6A4::::5.58:C|CP1A1:::sub::D;FMO1:::sub::D;CP3A4:::sub::D;CP2D6:::inh::D;CP2CJ:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;CP1A2:::sub::D||
Vildagliptin|ok_inv|DPP4:::inh:9.24:DC;DPP9::::7.18:C;DPP8::::6.09:C;SEPR::::5.43:C|||
Voglibose|inv|LYAG::::7.15:C;SUIS::RAT::7.15:C;LYAG::RAT::6.96:C;MGA:::inh:5.89:DC|||
Enoximone|ok_inv|BLM::::8.89:C;NFKB1::::6.1:C;PDE4A::::5.57:C;TSHR::::5.5:C;PDE3A:::inh:5.42:DC;CP3A4::::5.3:C;HCD2::::5.2:C|||
Dapoxetine|inv|5HT2C;5HT1B;5HT1A|CP2D6:::inh::D;CP3A4:::inh::D||
Cilansetron|inv|5HT3A::RAT::9.72:C;SGMR1::RAT::6.47:C;ACM1::RAT::6.04:C;5HT4R::RAT::6.02:C;5HT2C::RAT::5.31:C;CAC1C::RAT::5.27:C;HRH1::RAT::5.19:C;5HT2B::RAT::5.11:C;OPRM::RAT::5.07:C;5HT3A|||
Bepotastine|ok|HRH1:::ant::D|||
Vapreotide|exp_inv|SSR2:::ind::D;SSR5:::ago::D;NK1R:::ant::D|CP3A4:::inh::D||
Pegaptanib|ok_inv|NRP1|||
Milnacipran|ok_inv|SC6A4:::inh:8.19:DC;SC6A4::RAT::7.57:C;SC6A2:::inh:7.39:DC;NMDA:::inh::D|CP3A4:::inh::D||
Lucinactant|ok_inv||||
Ximelagatran|ok_out|THRB:::inh::D|CP2C9:::sub::D||
Nesiritide|ok_inv|ANPRA:::bin::D;ANPRB;ANPRC|||
Sitimagene_ceradenovec|inv||||
Flibanserin|ok_inv|5HT1A::RAT::7.93:C;5HT1A:::ago:6.2:DC;DRD4:::duo::D;5HT2A:::ant::D|CP3A4:::sub::D||
Oritavancin|ok_inv||CP3A4:::ind::D;CP2D6:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D||
Ceftobiprole|ok_inv|FTSI::ECOLI:::D;PBPX::STRPN:::D;MecA::STAAU:::D|||
Clevidipine|ok_inv|CAC1C::CAVPO::8.15:C;CAC1C;CAC1D;CAC1S;CAC1F|CHLE:::sub::D;CP3A4:::duo::D;CP2CJ:::inh::D;CP2E1:::sub::D;CP2D6:::sub::D;CP2C9:::inh::D||
rhThrombin|ok_inv||||
Itopride|inv|DRD2;ACES:::inh::D|||
Permethrin|ok_inv|TYDP1::::5.25:C;NR1I2;ESR1;SCN1A:::inh::D|CP2B6:::sub_ind::D||
Afamelanotide|ok_inv|MSHR::MOUSE::10.85:C;MC4R::::10.77:C;MSHR:::ago:10.64:DC;MC5R::MOUSE::10.52:C;MC3R::MOUSE::10.2:C;MC4R::MOUSE::10.01:C;MC3R::RAT::10.:C;MC3R::::9.89:C;MC5R::::9.64:C;ADA::::7.8:C|||
Defibrotide|ok_inv|AA1R;AA2AR;AA2BR|||
Ospemifene|ok_inv|ESR1:::duo::D|CP2D6:::inh::D;CP2B6:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D||
Crofelemer|ok|CFTR:::ant::D;ANO1:::ant::D|||
Acadesine|inv||||
Hemoglobin|ok_exp_inv||||
Iloperidone|ok|ADA2A::RAT::9.4:C;5HT2B::RAT::8.05:C;5HT2A::BOVIN::8.05:C;SGMR1::::7.19:C;DRD2::RAT::6.96:C;DRD2:::ant:6.96:DC;5HT1A::MOUSE::6.68:C;DRD1::MOUSE::6.12:C;ADA2C:::ant::D;HRH1:::ant::D;ADA1A:::ant::D;5HT7R:::ant::D;5HT6R:::ant::D;5HT1A:::ant::D;DRD4:::ant::D;DRD3:::ant::D;DRD1:::ant::D;5HT2A:::ant::D|CP2E1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D||
Lofexidine|ok_inv|ADA2C::::8.86:C;ADA2C::RAT::8.6:C;ADA2A:::ago:8.36:DC;NISCH::RAT::8.25:C;ADA2B::::7.17:C;5HT1A:::ago:6.9:DC;ADA1B::RAT::6.18:C;5HT1D:::ago::D;5HT2C:::ago::D;5HT7R:::ago::D;ADA1A:::ago::D|CP2CJ:::sub::D;CP1A2:::sub::D;CP2D6:::sub::D|S47A1:::inh::D;ABCB5:::inh::D|
Pirfenidone|ok_inv|BLM::::7.15:C;FURIN|CP1A2:::inh::D||
Ezogabine|ok_inv|KCNQ2::::6.37:DC;KCNQ2::MOUSE::5.89:C;KCNQ5;KCNQ4;KCNQ3|ARY2:::sub::D;UD19:::sub::D;UD14:::sub::D;UD13:::sub::D;UD11:::sub::D||
Afelimomab|inv|TNFA|||
Plitidepsin|inv||CP3A4:::sub::D;CP2A6:::sub::D;CP2E1:::sub::D;CP4AB:::sub::D||
Satraplatin|inv|DNA|||
Ingenol_mebutate|ok|KPCD:::lig:8.39:DC;KPCA:::lig::D|||
Belinostat|ok_inv|HDAC1,HDA10,HDA11,HDAC2,HDAC3,HDAC4,HDAC5,HDAC6,HDAC7,HDAC8,HDAC9:::inh:9.07,7.23,7.57,9.07,8.82,7.82,7.6,8.8,7.29,7.66,7.62:DC;HDAC1::::9.07:C;HDAC2::::9.07:C;HDAC3::::8.82:C;HDAC6::::8.8:C;HDAC4::::7.82:C;HDAC8::::7.66:C;HDAC9::::7.62:C;HDAC5::::7.6:C;HDA11::::7.57:C;HDAC7::::7.29:C;HDA10::::7.23:C|CP1A2:::ind::D;CP2C9:::inh::D;CP2C8:::inh::D;UD14:::inh::D|MDR1:::sub::D|
Ataluren|ok_inv|RORG::MOUSE::6.15:C|SO1B3:::inh::D;S22A8:::inh::D;S22A6:::inh::D;UD19:::sub::D||
Migalastat|ok_inv|AGAL::COFAR::8.52:C;AGAL::::7.15:DC;LYAG::::7.08:C;SUIS::::6.59:C;GLCM::::5.85:C;MGA::::5.82:C;AGALC::ASPNG::5.74:C;GDE::::5.:C|UD11:::sub::D||
Indacaterol|ok|ADRB2:::ago:8.82:DC;ADRB2::CAVPO::8.1:C;ADRB1::::7.04:C;DRD3::::5.98:C|UD11:::sub::D;CP3A4:::sub::D|MDR1:::sub::D|
Erdosteine|ok_inv||ADA:::inh::D||
Abaloparatide|ok_inv|PTH1R:::lig::D|||
Ancrod|ok_inv|FIBA|||
Pleconaril|inv|NR1I2::::6.6:C;CP2D6::::5.9:C;CP3A4::::5.2:C;Genome_polyprotein::9ENTO:::D|||
Trabectedin|ok_inv|DNA:::bin::D|PGH1:::sub::D;CP2CJ:::sub::D;CP2E1:::sub::D;CP2D6:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D||
Pretomanid|ok|INHA::MYCTU:::D;A0A0T9AZ62,A0A1K3GRG2,A0A045KKX4,A0A045ISQ8;LSR2::MYCTU:::D;EFPA::MYCTU:::D;Probable_fatty_acid_synthase_Fas_Fatty_acid_synthetase::MYCTU:::D|DDN::MYCTU:sub::D;CP3A4:::sub::D|S22A8:::inh::D|
Vintafolide|inv|FOLR2;FOLR3;FOLR1|||
Crisaborole|ok_inv|PDE4A:::inh:6.96:DC;PDE7A::::6.14:C;PDE1A::::5.21:C;PDE3A::::5.19:C;PDE4D:::inh::D;PDE4C:::inh::D;PDE4B:::inh::D|CP2C9:::inh::D;CP2C8:::inh::D;CP2B6:::inh::D||
Beraprost|inv|PI2R|CP2C8:::sub::D||
Cobimetinib|ok_inv|MP2K1:::inh:9.05:DC|MDR1:::sub::D;CP3A4:::sub::D|ABCG2:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D|
Silver_sulfadiazine|ok_vet|DNA:::bin::D|||
Methsuximide|ok|CAC1G:::inh::D|CP2CJ:::inh::D||
Fibrinolysin|inv|PAI1;UROK|||
Glatiramer|ok_inv|2B11:::bin::D|||
Gallium_nitrate|ok_inv|RIR2:::inh::D;VATB2:::inh::D;OSTCN:::ant::D;Hydroxylapatite:::mod::D;Protein_tyrosine_phosphatase::9GAMM:inh::D;IL1B:::ant::D||TFR1|TRFE:::sub::D
Ibudilast|inv|BLM::::7.6:C;CP2D6::::7.4:C;PDE4A:::inh:7.27:DC;PDE4B:::inh:7.19:DC;PDE4D:::inh:6.78:DC;PDE4C:::inh:6.62:DC;CP1A2::::6.2:C;CP2CJ::::5.5:C;CP3A4::::5.1:C;PDE3A:::inh::D|||
Rotigotine|ok|DRD2:::ago:10.22:DC;DRD3:::ago:8.4:DC;DRD2::BOVIN::7.82:C;DRD1:::ago:7.55:DC;DRD4:::ago:7.26:DC;DRD1::BOVIN::6.3:C;ADA2B:::ant::D;5HT1A:::ago::D;DRD5:::ago::D|CP2D6:::inh::D;CP3A4:::sub::D||
Samarium_153Sm_lexidronam|ok_inv||||
Hepatitis_B_Immune_Globulin|ok_inv|HBsAg::HBV:::D|||
Vandetanib|ok|RIPK2::::8.34:C;EGFR:::inh:8.32:DC;EGFR:G719S::inh:8.23:DC;VGFR2::::8.2:C;EGFR:L858R::inh:8.06:DC;ABL1:Y253F:::8.05:C;EGFR:G719C::inh:8.02:DC;ABL1:H396P:::8.01:C;EGFR:L861Q::inh:7.96:DC;DDR1::::7.96:C;ABL1:E255K:::7.89:C;RET:M918T:::7.85:DC;ABL1:M351T:::7.82:C;ABL1:Q252H:::7.8:C;ABL1::::7.8:C;LCK::::7.77:C;ABL1:T315I:::7.7:C;RET::::7.7:DC;VGFR1::::7.66:C;PTK6:::inh:7.48:DC;ABL1:F317L:::7.48:C;KIT:A829P:::7.47:C;SRC::::7.36:C;MP2K5::::7.31:C;EPHA6::::7.3:C;STK35::::7.25:C;TYRO3::::7.2:C;BLK::::7.18:C;ABL2::::7.16:C;IRAK4::::7.12:C;EPHB6::::7.12:C;STK10::::7.09:C;GAK::::7.07:C;PGFRB::::7.06:C;EPHA8::::7.04:C;SLK::::7.02:C;EGFR:T790M::inh:7.:DC;ROCK2::::7.:C;LYN::::6.96:C;YES::::6.92:C;KIT:L576P:::6.85:C;ACVR1::::6.82:C;M4K4::::6.8:C;ERBB3::::6.8:C;PGFRA::::6.8:C;FRK::::6.77:C;ABL1:F317I:::6.77:C;KIT:V559D:::6.74:C;FLT3:K663Q:::6.72:C;EPHA1::::6.64:C;EGFR:L858R-T790M::inh:6.64:DC;VGFR3::::6.63:C;EPHA5::::6.62:C;FGFR3::::6.62:C;KS6A6::::6.62:C;BMR1B::::6.62:C;UFO::::6.6:C;KIT::::6.59:C;FGR::::6.57:C;KIT:D816V:::6.54:C;EPHB1::::6.54:C;M4K5::::6.5:C;DDR2::::6.49:C;MKNK1::::6.44:C;HCK::::6.44:C;FYN::::6.44:C;KS6A1::::6.4:C;LTK::::6.4:C;KIT:D816H:::6.38:C;SIK2::::6.37:C;EPHB2::::6.36:C;ACVL1::::6.33:C;ERBB4::::6.32:C;TBA1A::RAT::6.32:C;EPHB4::::6.28:C;KIT:V559D-V654A:::6.25:C;FGFR1::::6.25:C;FLT3:D835H:::6.25:C;TIE2:::inh:6.25:DC;RIPK4::::6.21:C;PLK4::::6.21:C;FLT3:D835Y:::6.08:C;FLT3::::6.07:C;M3K19::::6.01:C;MP2K1::::6.:C;FGFR2::::5.96:C;MP2K2::::5.96:C;EPHA2::::5.96:C;PHKG1::::5.96:C;CSF1R::::5.92:C;IRAK1::::5.92:C;FLT3:N841I:::5.92:C;BTK::::5.9:C;FLT3:R834Q:::5.89:C;MERTK::::5.85:C;STK33::::5.85:C;MK06::::5.82:C;TIE1::::5.82:C;AURKC::::5.82:C;KC1E::::5.82:C;M4K3::::5.82:C;EPHA4::::5.8:C;M4K2::::5.8:C;KS6B1::::5.8:C;ALK::::5.8:C;MKNK2::::5.77:C;COQ8B::::5.77:C;CTRO::::5.74:C;EPHA3::::5.74:C;SRMS::::5.72:C;SIK1::::5.72:C;KIT:V559D-T670I:::5.7:C;LRRK2::::5.7:C;MRCKG::::5.66:C;TNIK::::5.64:C;FGFR4::::5.64:C;EPHA7::::5.62:C;AURKB::::5.6:C;MK14::::5.6:C;CSK::::5.6:C;MRCKB::::5.6:C;MRCKA::::5.59:C;ERBB2::::5.59:C;TNI3K::::5.55:C;AAPK1::::5.52:C;M3K4::::5.52:C;MINK1::::5.47:C;RON::::5.47:C;TESK1::::5.43:C;TXK::::5.43:C;SIK3::::5.41:C;MET:Y1235D:::5.39:C;CDK7::::5.39:C;HUNK::::5.39:C;COQ8A::::5.35:C;ST32A::::5.3:C;M3K20::::5.29:C;M4K1::::5.26:C;MET::::5.24:C;ULK3::::5.19:C;FGFR3:G697C:::5.16:C;PHKG2::::5.1:C;VEGFA:::inh::D|CP3A4:::sub::D;FMO3:::sub::D;FMO1:::sub::D|S22A2:::inh::D;ABCG2:::inh::D;MRP1:::inh::D|ALBU:::bin::D;A1AG1:::bin::D
keyhole_limpet_hemocyanin|ok_inv|IL2|||
Ecallantide|ok_inv|KLKB1:::inh::D|||
Pimavanserin|ok_inv|5HT2A:::ANT::D;DRD2|||
Romiplostim|ok|TPOR:::ago::D|||
Obiltoxaximab|ok||||
Dexlansoprazole|ok_inv|TAU::::8.6:C;ACM1::RAT::7.25:C;TSHR::::6.9:C;LMNA::::6.9:C;ATP4A:::inh:6.4:DC;PHOP1::::6.36:C;HCD2::::6.3:C;NPC1::::5.64:C;RAB9A::::5.64:C;CP2D6::::5.54:C;AGAL::::5.3:C;FAS::::5.28:C;CP2C8::::5.24:C;CP1A2::::5.19:C;HIF1A::::5.1:C;I23O2::MOUSE::5.09:C;DDAH1;ATP4B:::inh::D|CP2CJ:::inh:7.:DC;CP3A4:::sub::D||
Ragweed_pollen_extract|ok_inv||||
Histamine|ok_inv|HRH3::CAVPO::9.84:C;HRH1::CAVPO::9.11:C;HRH4:::ago:8.8:DC;HRH3:::ago:8.39:DC;HRH3::RAT::8.2:C;HRH1::RAT::8.:C;HRH1:::ago:7.89:DC;HRH4::MOUSE::7.38:C;HRH4::RAT::7.2:C;HRH3::MOUSE::7.17:C;HRH2:::ago:6.33:DC;LMNA::::6.05:C;HRH2::CAVPO::6.:C;FFP::BACIU::5.:C;VMAT2|HNMT:::sub::D|S22A5:::inh::D;S22A3:::inh::D;S22A1;S22A2:::inh::D|
Iodine|ok_inv|NU5M|||
Carbopol_974P|ok_inv||||
Tetrachlorodecaoxide|ok_inv|MAEA;C163A|||
Corticorelin|inv||DOPO:::ind::D||
Albinterferon_Alfa_2B|inv||CP1A2:::inh::D||
Briakinumab|inv|IL12B;IL23A|||
Telaprevir|ok_out|CMA1::::7.59:C;CELA1::::7.52:C;CATB::::6.68:C;CATS::::6.52:C;CATK::::6.2:C;ELNE::::6.17:C;CATL2::::5.87:C;CATL1::::5.46:C;PLMN::::5.06:C;SO2B1:::inh::D;SO1B1:::inh::D;Genome_polyprotein::9HEPC:inh::D|CP3A4:::inh::D|MDR1:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Mipomersen|ok_inv|mRNA:::bin::D|||
Brivaracetam|ok_inv|SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A,SCN1B,SCN2B,SCN3B,SCN4B:::inh::D;SV2A|CP2C9:::sub::D;CP2B6:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D||
Ramucirumab|ok_inv|VGFR2:::ant::D|||
Sodium_stibogluconate|ok_inv|TOP1:::inh::D|||
Apremilast|ok_inv|PDE4A::::7.13:C;Phosphodiesterase_isozyme_4:::ant::D|CP1A2:::sub::D;CP2A6:::sub::D;CP3A4:::sub::D|MDR1:::sub::D|
Ustekinumab|ok_inv|IL12B:::inh::D;IL12B:::inh::D|||
Trastuzumab_emtansine|ok_inv|ERBB2:::abo::D|CP3A4:::inh::D;CP3A5:::sub::D|MDR1:::sub::D|
Thrombomodulin_Alfa|ok_inv|THRB:::inh::D;FA5|||
Perflubron|inv|LMNA::::6.15:C|||
Serelaxin|inv||||
Abiraterone|ok|CP17A:::inh:8.54:DC;CP17A::RAT::7.9:C;C11B1::::5.79:C;C11B2::::5.76:C|CP3A4:::inh:5.57:DC;CP2C9:::inh::D;CP2CJ:::inh::D;CP1A2:::inh::D;CP2C8:::inh::D;CP2D6:::inh::D;ST2A1:::sub::D|MRP1:::inh::D|A1AG1:::bin::D;ALBU:::bin::D
Parathyroid_hormone|ok_inv|PTH1R:::act::D;PTH2R:::act::D|||
Inotuzumab_ozogamicin|ok_inv|CD22:::abo::D||MDR1:::sub::D|
Obeticholic_acid|ok|NR1H4:::ago:7.07:DC;GPBAR::::7.:C|CP1A2:::inh::D;BAAT:::sub::D||
Eteplirsen|ok_inv|DMD:::bin::D|||
Cariprazine|ok_inv|DRD3:::ago:10.02:DC;DRD2:::ago:9.39:DC;5HT1A:::ago:8.51:DC;5HT2A:::ant:7.66:DC;DRD4::::6.96:C;DRD1::::5.68:C;HRH1:::ant::D;5HT2B:::ant::D|CP2D6:::sub::D;CP3A4:::sub::D||
Olaratumab|ok_inv|PGFRA:::ant::D|||
Lumateperone|ok_inv|5HT2A:::ant::D;DRD2:::pag::D;DRD1;SC6A4:::inh::D;NMDE2|AKCL2;CP3A4;CP2C8;CP1A2;UD11;UD14;UDB15;AK1C1;AK1BA;AK1C4||
Caplacizumab|ok_inv|VWF|||
Cenobamate|ok_inv||UD2B7:::sub::D;UD2B4:::sub::D;CP2E1:::sub::D;CP2A6:::sub::D;CP2B6:::duo::D;CP2CJ:::inh::D;CP3A4:::duo::D;CP3A5:::inh::D;CP2C8:::ind::D||ALBU:::bin::D
Sertindole|ok_out|5HT2C:::ant:9.7:DC;5HT2A::RAT::9.7:C;ADA1B::MESAU::9.48:C;ADA1A::BOVIN::9.43:C;5HT2B::RAT::9.41:C;DRD2:::ant:9.35:DC;DRD2::RAT::9.35:C;HRH1::::9.29:C;5HT2C::RAT::9.29:C;5HT2A:::ant:9.22:DC;ADA1D::RAT::9.18:C;ADA1B::RAT::8.85:C;ADA1A::::8.74:DC;DRD3::::8.59:C;KCNH2:::inh:8.57:DC;ADA1A::RAT::8.47:C;5HT6R:::ant:8.3:DC;DRD4::::7.96:C;DRD1::RAT::7.92:C;5HT1A::::7.48:C;5HT1B::::7.25:C;DRD1::::6.68:C;ADA2A::::5.77:C;KCNA5::::5.7:C;SCN1A::::5.64:C;CAC1C::::5.2:C;MDR1::::5.19:C;ADA1D;ADA1B|CP3A4:::sub::D;CP2D6:::sub::D||
Spiramycin|ok|RL3::STRP1:ant::D|||
Sulfathiazole|ok_vet|DHPS::ECOLI::5.6:C;Dihydropteroate_synthetase::PLAFA:inh::D|CP19A:::ind::D||
Mianserin|ok_inv|ADA1A::RAT::10.15:C;HRH1:::ant:9.76:DC;5HT2A:::ant:9.3:DC;5HT2C:::ant:9.22:DC;HRH1::CAVPO::9.07:C;5HT2B::RAT::8.96:C;5HT2C::RAT::8.85:C;5HT2A::RAT::8.82:C;ADA2C:::ant:8.42:DC;5HT2B:::bin:8.33:DC;ADA2A:::ant:8.32:DC;ADA2A::BOVIN::7.77:C;ADA2B:::ant:7.62:DC;ADA1B::RAT::7.55:C;5HT6R:::bin:7.4:DC;ADA1D::::7.39:C;ADA1A::BOVIN::7.37:C;ADA2C::RAT::7.27:C;5HT7R:::ant:7.25:DC;5HT7R::RAT::7.2:C;5HT3A::RAT::7.15:C;LMNA::::6.8:C;SC6A2:::inh:6.79:DC;ACM5::::6.64:C;FFP::BACIU::6.63:C;ADA1A,ADA1B,ADA1D:::ant:6.6,,7.39:DC;ADA1A::::6.6:C;5HT3B::MOUSE::6.6:C;DRD1,DRD5:::bin:6.57,:DC;DRD1::::6.57:C;ACM4::::6.54:C;ACM3::::6.53:C;ACM1::::6.46:C;ACM2::::6.42:C;5HT1D::::6.42:C;5HT1A:::inh:6.4:DC;5HT1A::RAT::6.3:C;5HT1B::RAT::6.24:C;DRD2::RAT::6.08:C;HRH2::CAVPO::6.06:C;HRH2::::6.:C;SC6A4:::inh:5.96:DC;5HT3A::::5.85:C;DRD1::RAT::5.85:C;DRD3::RAT::5.82:C;ACM5::RAT::5.72:C;DRD2:::ant:5.66:DC;DRD3:::bin:5.55:DC;SC6A4::RAT::5.54:C;DRD4::::5.48:C;SCN1A::::5.26:C;SC6A3:::bin::D;OPRK:::ago::D;5HT1F:::bin::D;HRH4:::bin::D|CP2B6:::sub::D;CP1A2:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D||
Teicoplanin|ok_inv|D::G+Bac:inh::D|||
Sulfadimethoxine|ok_vet|LMNA::::8.74:C;LEF::BACAN::6.6:C;5HT6R::::6.21:C;CYSP::TRYCR::5.2:C|CP2C9:::inh::D||
Acetylcysteine|ok_inv|THB::::6.25:C;BLM::::6.:C;RECQ1::::5.85:C;NFKB1::::5.35:C;NMD3A:::act::D;NMDE4:::act::D;NMDE1:::act::D;NMDZ1:::act::D;NMDE2:::act::D;IKKA:::inh::D;IKKB:::inh::D;ACY1:::lig::D;NAPQI:::reducer::D;XCT:::act::D;GSHB:::sti::D||S22A6;SO1B1:::inh::D|
Nylidrin|ok|INAR2:::ago::D;CAC1I:::duo::D|CP3A4:::sub::D;COMT:::ind::D||
Pizotifen|ok|5HT2C:::ant:8.85:DC;ACM1:::ant:8.7:DC;5HT2B:::ant:8.7:DC;DRD2::::8.62:C;5HT2A:::ant:8.12:DC;5HT7R::::7.6:C;ADA2C:::ant::D;ADA2B:::ant::D;ADA2A:::ant::D;ADA1D:::ant::D;ADA1B:::ant::D;ADA1A:::ant::D;HRH1:::ant::D;5HT1D:::ant::D;5HT1B:::ant::D;5HT1A:::ant::D;ACM3:::ant::D;ACM2:::ant::D|UDB10:::sub::D||
Pentaerythritol_tetranitrate|ok|AL1A1::::5.8:C;Free_radicals:::ant::D;HBB:::ago::D;HBA:::ago::D|ALDH2:::sub::D;NOS3:::ind::D;GCYA2:::ind::D||
Rimonabant|ok_inv|CNR1:::ant:9.96:DC;CNR1::RAT::9.77:C;CNR2::::8.96:C;CNR1::MOUSE::8.82:C;CP2C9::::8.28:C;CNR2::MOUSE::6.43:C;MRP1::::5.85:C;GPR55::::5.7:DC;KCNH2::::5.55:C;MRP4::::5.4:C;GPR18::::5.:C|CP3A4:::sub::D||
Garenoxacin|inv||CP1A2:::inh::D||
Canakinumab|ok_inv|IL1B:::bin::D|||
Noscapine|ok_inv|CP2CJ::::6.8:C;TBB4B::::5.73:C;S22A2::::5.59:C;SGMR1|CP2C9:::inh:6.9:DC;CP3A4:::inh:5.7:DC||
Romidepsin|ok_inv|HDAC1:::ant:9.7:DC;HDAC2:::ant:9.:DC;HDAC3::::8.52:C;HDAC6:::inh:6.7:DC;HDAC4:::inh:6.29:DC;MRP1|CP2CJ:::sub::D;CP2B6:::sub::D;CP1A1:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|SO1B3:::sub::D;MDR1:::sub::D|
Ipilimumab|ok|CTLA4|||
Pixantrone|ok_inv||||
Icatibant|ok_inv|BKRB2:::ant:10.6:DC;BKRB2::RAT::10.11:C;BKRB2::CAVPO::10.05:C;AMPN:::inh::D|||
Tedisamil|inv|KCNH2::::5.6:C|||
Rufinamide|ok|SCN9A:::mod::D;GRM5:::inh::D|CP3A4:::sub_ind::D;CP2E1:::inh::D;EST1:::sub::D||ALBU:::sub::D
Lasofoxifene|ok_inv|ESR2:::ago:10.:DC;ESR1:::ant:8.89:DC;ESR1::RAT::7.95:C;CNR2:::ANT::D|||
Alogliptin|ok|DPP4:::inh:9.:DC|CP2D6:::sub::D;CP3A4:::sub::D||
Tapentadol|ok|OPRM:::ago:6.8:DC;SC6A4:::inh::D;5HT3A;OPRD;OPRK;SC6A2:::inh::D|CP2CJ:::sub::D;CP2C9:::sub::D;CP2D6:::inh::D;UD2B7:::sub::D;UD19:::sub::D||
Vorhyaluronidase_alfa|ok_inv|Hyaluronan;TGFB1:::inh::D|||ALBU:::inh::D
Sugammadex|ok||||
Silodosin|ok|ADA1A:::ant:10.44:DC;ADA1A::RAT::9.1:C;ADA1D:::ant:8.7:DC;ADA1B:::ant:7.7:DC;ADA1B::RAT::7.05:C;KCNH2::::5.1:C|UD2B7:::sub::D;CP3A4:::sub::D|MDR3:::sub::D;MDR1:::sub::D|
Prasugrel|ok|P2Y12:::ant::D|CP2CJ:::sub::D;CP2C9:::sub::D;CP2B6:::sub::D;CP3A4:::sub::D;EST2:::sub::D||ALBU:::sub::D
Eltrombopag|ok|TPOR:::ago:7.42:DC;KCNH2::::6.2:C;SO2B1::::5.07:C|UD19:::inh::D;UD13:::sub::D;UD11:::inh::D;CP1A2:::sub::D;CP2C8:::inh::D|ABCG2:::inh::D;SO1B1:::inh::D|
Doripenem|ok_inv|CAC1C::::5.7:C;Penicillin_binding_protein_4::STAAU:ant::D;Cell_division_protein::PSEAI:ant::D;MRDA::ECOLI:ant::D;PBPB::ECOLI:ant::D;PBPA::ECOLI:ant::D|DPEP1:::sub::D|S22A8:::sub::D|
Tolvaptan|ok|V2R:::ant:9.37:DC;V1AR:::ant::D|CP3A4:::sub::D|MDR1:::inh::D|
Regadenoson|ok_inv|AA2AR:::ago:6.54:DC;AA2AR::RAT::6.54:C;AA1R::::5.42:C;AA3R::::5.:C;AA2BR::::5.:C|||
Ferumoxytol|ok_inv|||TRFE:::tra::D;FRIL:::sto::D;FRIH:::sto::D|
Asenapine|ok|5HT1A:::ant::D;5HT1B:::ant::D;5HT2A:::ant::D;5HT2B:::ant::D;5HT2C:::ant::D;5HT5A:::ant::D;5HT6R:::ant::D;5HT7R:::ant::D;DRD2:::ant::D;DRD3:::ant::D;DRD4:::ant::D;DRD1:::ant::D;ADA1A:::ant::D;ADA2A:::ant::D;ADA2B:::ant::D;ADA2C:::ant::D;HRH1:::ant::D;HRH2:::ant::D;ADRB1:::ant::D;ADRB2:::ant::D|UD14:::sub::D;CP1A2:::sub::D;CP2D6:::inh::D;CP3A4:::sub::D||ALBU:::bin::D;A1AG1:::bin::D
Vernakalant|ok_inv|SCN5A:::inh::D;KCNA5:::inh::D;KCND3:::inh::D;KCNH2:::inh::D|CP2D6:::inh::D||
Lacosamide|ok|SCN9A::::6.74:DC;CAH2::::6.48:C;CAH5B::::6.47:C;CAH9::::6.45:C;CAH1::::6.44:C;CAH3::::6.43:C;CAH6::::6.39:C;SCN3A::RAT::6.38:C;CAH15::MOUSE::6.34:C;CAH14::::6.33:C;CAH4::::6.28:C;CAH13::::5.92:C;CAH12::::5.43:C;CAH7::::5.35:C;CAH5A::::5.34:C;SCNAA;SCN3A|CP3A4:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D||
Dalbavancin|ok_inv|D::G+Bac:bin::D|||
Rivaroxaban|ok|FA10:::ant:9.4:DC;FA10::RABIT::6.29:C;ST14::::5.47:C|CP3A5:::sub::D;CP2J2:::sub::D;CP3A4:::sub::D|ABCG2:::sub::D;MDR1:::sub::D|
Nalmefene|ok_out|OPRK:::pag:10.08:DC;OPRM:::ant:9.62:DC;OPRM::RAT::9.54:C;OPRD:::ant:9.04:DC;OPRK::CAVPO::8.7:C;OPRD::RAT::8.47:C|UD18:::sub::D;UD13:::sub::D;UD2B7:::sub::D||
Ridaforolimus|inv|MTOR|CP3A4:::inh::D||
Maribavir|inv|UL97::HCMVT:::D;UL97::HCMVA:::D|||
Avanafil|ok|PDE5A::CANLF::8.28:C;PDE5A:::inh:8.16:DC|CP3A4:::sub::D||
Eflornithine|ok_out|DCOR:::ant::D|||
Arzoxifene|ok_inv|ESR1::::9.7:DC;ESR2::::7.18:DC|||
Hexaminolevulinate|ok||||
Droxidopa|ok_inv|NR1I2::::8.4:C;PH4H:::inh::D;ADRB3:::ago::D;ADRB2:::ago::D;ADRB1:::ago::D;ADA2C:::ago::D;ADA2B:::ago::D;ADA2A:::ago::D;ADA1D:::ago::D;ADA1B:::ago::D;ADA1A:::ago::D|DDC:::sub::D|MOT10:::inh::D;SC6A2:::sub::D|
Amrubicin|inv|TOP2A;DNA|NCPR:::sub::D;CBR1:::sub::D|ABCB5:::sub::D|
Tolperisone|inv|SGMR1::::8.25:C;ADA2B::::6.34:C|CP1A2:::sub::D||
Lonidamine|inv|AMPC::ECOLI::6.25:C;CP3A4::::5.6:C;NPSR1::::5.5:C;HXK1;CFTR|||
Udenafil|ok_inv|PDE5A:::inh::D|CP3A4:::sub::D;CP3A5:::sub::D||
Sitaxentan|ok_out|EDNRA:::ant:9.37:DC;EDNRA::RAT::9.37:C;EDNRB:::ant:8.01:DC|CP2CJ:::inh::D;CP3A4:::inh::D;CP2C9:::inh::D||
Sulodexide|ok_inv|HEP2:::ago::D;ANT3:::pot::D|||
Tocilizumab|ok|IL6RA:::abo::D|CP3A4:::ind::D||
Alvimopan|ok_inv|OPRM:::ant:9.33:DC;OPRD:::ant:7.92:DC;OPRK:::ant:7.:DC;CAC1C::::5.3:C|||
Levocetirizine|ok|HRH1:::ant::D|CP3A4:::sub::D|S22AB:::sub::D|ALBU:::bin::D
Ziconotide|ok|CAC1B::::6.3:C|CP3A4:::sub::D||
Teriparatide|ok_inv|PTH1R:::bin:9.52:DC|||
Temsirolimus|ok|MTOR:::inh:5.75:DC|CP2D6:::inh::D;CP3A7:::sub::D;CP3A5:::inh::D;CP3A4:::sub::D|MDR1:::inh::D|
Amisulpride|ok_inv|DRD2:::ant:8.52:DC;DRD3:::ant:8.4:DC;5HT7R:::ant:7.6:DC;ADA2C::RAT::6.9:C;5HT2B::::6.5:C;5HT2A:::ant:6.2:DC;LMNA::::5.4:C|||
Simeprevir|ok|CATS::::6.1:C;NS3_protease::9HEPC:inh::D|CP3A4:::inh::D;CP1A2:::inh::D|ABCBB:::inh::D;NTCP:::inh::D;SO2B1:::sub::D;ABCG2:::inh::D;MRP2:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;MDR1:::inh::D|ALBU:::bin::D
Dapagliflozin|ok|SC5A2:::ant:9.31:DC;SC5A4::::8.87:C;SC5A2::RAT::8.52:C;SC5A1::::8.49:C;SC5AB::::6.42:C|UD2B7:::sub::D;UD2B4:::sub::D;UD19:::sub::D;CP3A4:::sub::D;CP2D6:::sub::D;CP2C9:::sub::D;CP2A6:::sub::D;CP1A2:::sub::D;CP1A1:::sub::D|MDR1:::sub::D|
Motavizumab|inv||||
Elotuzumab|ok|SLAF7:::mod::D|||
Saxagliptin|ok|DPP4:::inh:9.22:DC;DPP9::::7.15:C;DPP8::::6.89:C|CP3A5:::sub::D;CP3A4:::sub::D|S22A8:::sub::D;SO4C1:::sub::D;MRP1:::sub::D|
Iclaprim|inv|DYR::STAAU::10.1:C;DYR::::8.1:DC;DYR::PNECA::5.62:C|||
rsPSMA_Vaccine|ok_inv||||
Pertuzumab|ok|ERBB2:::abo::D|||
Rilonacept|ok_inv|IL1B:::bin::D;IL1A:::bin::D;IL1RA:::bin::D|||
Xaliproden|inv|5HT1A|||
Bazedoxifene|ok_inv|ESR1:::duo:9.22:DC;ESR2::::8.42:DC|UD110:::sub::D;UD18:::sub::D;UD14:::sub::D||
Telavancin|ok||||
Ambrisentan|ok_inv|EDNRA:::ant:7.66:DC;EDNRA::RAT::7.09:C;EDNRB:::ant:5.92:DC|CP3A5:::sub::D;UD13:::sub::D;UD2B7:::sub::D;UD19:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D|SO1B3:::sub::D;SO1B1:::sub::D;MDR1:::sub::D|
Human_C1_esterase_inhibitor|ok|C1R:::inh::D;C1S:::inh::D;KLKB1:::inh::D;FA12:::inh::D;THRB:::inh::D;FA11:::inh::D;TPA:::inh::D|||
Doxercalciferol|ok|VDR:::sup::D|CP27A:::act::D||
Oxymetholone|ok_ill|AL1A1::::7.15:C;ANDR::RAT::6.86:C;LEF::BACAN::5.4:C;NPSR1::::5.2:C;RORG::MOUSE::5.:C;ANFB;ANDR:::ago::D|CP343:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D;S5A1:::act::D;CP2D6:::inh::D;AOFA:::ind::D||SHBG;ALBU
Armodafinil|ok_inv|LMNA::::8.74:C;DRD2::::8.68:C;SC6A3:::ant:6.19:DC;SC6A3::RAT::5.6:C|CP2C9:::inh::D;CP2B6:::ind::D;CP1A2:::ind::D;CP3A5:::ind::D;CP3A4:::ind::D;CP2CJ:::inh::D||
Etravirine|ok|CYSP::TRYCR::5.4:C;MRP3::::5.29:C;ABCG2::::5.22:C;MRP2::::5.11:C;MRP1::::5.07:C;POL::HV1H2:::D;POL::HV1B1:::D|CP2CJ:::inh::D;CP2C9:::duo::D;CP3A4:::sub_ind::D|MDR1:::ind:5.12:DC;MDR3:::inh::D|
Calfactant|ok||||
Tyloxapol|ok_inv|LIPL:::inh::D|||
Cangrelor|ok|P2Y12:::inh:9.4:DC|||
Clomethiazole|inv|LMNA::::7.65:C;CP2C9::::5.6:C;GBRA1|CP2CJ:::sub:5.1:DC;CP3A4:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D||
Propentofylline|inv|LMNA::::7.3:C;NFKB1::::5.6:C;ACES::::5.19:C;PDE4A|CP1A2:::sub::D||
Prucalopride|ok|5HT4R:::ago:8.6:DC;5HT4R::RAT::7.59:C;5HT3A::::5.4:C|CP3A4:::sub::D|MDR1:::sub::D|ALBU:::bin::D
Etilevodopa|inv||||
Pazopanib|ok|KIT:L576P::inh:8.74:DC;PGFRB:::inh:8.7:DC;KIT:V559D::inh:8.64:DC;KIT:::inh:8.55:DC;VGFR2:::inh:8.5:DC;PGFRA:::inh:8.31:DC;KIT:V559D-T670I::inh:8.19:DC;CSF1R::::8.1:C;VGFR1:::inh:8.:DC;VGFR3::::7.57:DC;KIT:V559D-V654A::inh:7.52:DC;KIT:A829P::inh:7.48:DC;TAOK3::::7.35:C;DDR2::::7.3:C;DDR1::::7.24:C;RET::::7.1:C;EPHB6::::7.09:C;STK10::::7.08:C;FGFR1::::6.85:C;TTK::::6.82:C;GAK::::6.7:C;FGFR2::::6.68:C;SLK::::6.62:C;TAOK1::::6.62:C;RIPK1::::6.59:C;RET:M918T:::6.57:C;PI42C::::6.55:C;M3K9::::6.54:C;M3K2::::6.54:C;PLK4::::6.54:C;TNIK::::6.51:C;M4K4::::6.5:C;ABL1::::6.5:C;STK16::::6.44:C;CDPK1::PLAF7::6.43:C;ABL1:H396P:::6.42:C;LIMK2::::6.41:C;NEK2::::6.4:C;BRAF:V600E:::6.37:C;STK36::::6.33:C;ABL1:Y253F:::6.32:C;MP2K5::::6.32:C;KIT:D816V::inh:6.3:DC;MK08::::6.3:C;LCK::::6.3:C;ABL1:Q252H:::6.28:C;ABL1:M351T:::6.25:C;RIPK2::::6.24:C;MP2K4::::6.23:C;FGFR3:G697C::inh:6.21:DC;RIOK2::::6.21:C;AURKA::::6.2:C;TIE1::::6.15:C;BRAF::::6.14:C;LIMK1::::6.14:C;M3K11::::6.13:C;FGFR3:::inh:6.13:DC;FLT3:K663Q:::6.13:C;AURKC::::6.12:C;M4K1::::6.12:C;FRK::::6.12:C;ABL1:E255K:::6.1:C;IRAK3::::6.1:C;FLT3:D835Y:::6.09:C;RAF1::::6.05:C;LYN::::6.05:C;ROS1::::6.04:C;M3K19::::6.03:C;ACES::::6.03:C;PI4KB::::6.02:C;TNK1::::6.01:C;KIT:D816H::inh:6.:DC;BMR1B::::6.:C;FLT3::::5.96:C;FLT3:D835H:::5.96:C;CDK16::::5.92:C;AURKB::::5.9:C;CD11A::::5.89:C;FES::::5.85:C;MET::::5.8:C;M4K3::::5.8:C;FLT3:N841I:::5.8:C;FGR::::5.8:C;LTK::::5.8:C;ALK::::5.8:C;JAK2::::5.77:C;TAOK2::::5.74:C;MK10::::5.72:C;E2AK2::::5.72:C;PI51C::::5.72:C;IGF1R::::5.7:C;MK09::::5.7:C;MYLK2::::5.7:C;FYN::::5.7:C;M3K10::::5.68:C;CD11B::::5.68:C;MET:Y1235D:::5.68:C;KCC1A::::5.68:C;ABL1:T315I:::5.68:C;SIK1::::5.66:C;PTK6::::5.64:C;RET:V804M:::5.64:C;AVR2B::::5.62:C;SRMS::::5.6:C;TXK::::5.59:C;BLK::::5.59:C;FER::::5.57:C;M4K2::::5.57:C;ABL1:F317L:::5.57:C;SRC::::5.55:C;FGFR4::::5.55:C;AAK1::::5.54:C;M3K1::::5.54:C;M4K5::::5.52:C;TGFR2::::5.52:C;ABL2::::5.52:C;ACK1::::5.5:C;MERTK::::5.48:C;TIE2::::5.48:C;MET:M1250T:::5.47:C;TYK2::::5.47:C;KCC1G::::5.43:C;MARK3::::5.4:C;CDK7::::5.4:C;MP2K6::::5.39:C;NLK::::5.36:C;KSYK::::5.33:C;YES::::5.3:C;FAK1::::5.3:C;HCK::::5.24:C;IRAK1::::5.23:C;RET:V804L:::5.23:C;JAK3::::5.16:C;SIK2::::5.14:C;NEK5::::5.14:C;BMP2K::::5.06:C;FLT3:R834Q:::5.02:C;SH2B3:::inh::D;FGF1:::inh::D;ITK:::inh::D|CP1A2:::sub::D;CP2C8:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D|UD11:::inh::D;SO1B1:::inh::D;ABCG2:::sub::D;MDR1:::sub::D|
Ceftaroline_fosamil|ok_inv||||
Agomelatine|ok_inv|MTR1A:::ago:10.22:DC;MTR1B:::ago:10.:DC;MTR1C::CHICK::9.28:C;5HT2C:::ant:6.2:DC|CP2C9:::inh::D;CP1A2:::sub::D||
Midostaurin|ok_inv|FLT3:K663Q::ant:8.7:DC;FLT3:N841I::ant:8.22:DC;FLT3:D835H::ant:8.17:DC;KIT:D816V::ant:8.11:DC;EGFR:L858R-T790M:::8.06:C;PKN1::::8.03:C;TBK1::::8.03:C;EGFR:T790M:::8.01:C;FLT3:::ant:7.96:DC;JAK3::::7.92:C;FLT3:R834Q::ant:7.92:DC;M3K9::::7.82:C;PKN2::::7.82:C;M3K19::::7.82:C;FLT3:D835Y::ant:7.82:DC;KIT:D816H::ant:7.8:DC;STK4::::7.77:C;M3K11::::7.77:C;AURKA::::7.71:C;KCC2A::::7.7:C;RET:V804M:::7.7:C;MARK3::::7.68:C;RET:V804L:::7.57:C;KCC2D::::7.44:C;E2AK4::::7.41:C;STK3::::7.4:C;NUAK1::::7.39:C;KIT:L576P::ant:7.39:DC;SRPK1::::7.38:C;KIT:A829P::ant:7.37:DC;AAK1::::7.32:C;GRK7::::7.32:C;PRP4::::7.26:C;PRP4B::::7.26:C;AURKB::::7.21:C;NUAK2::::7.2:C;PLK4::::7.18:C;KKCC2::::7.14:C;KGP2::::7.13:C;SRPK3::::7.1:C;TNK1::::7.08:C;RK::::7.07:C;KSYK::::7.06:C;JAK2::::7.03:C;SIK3::::7.01:C;RIOK2::::7.01:C;DYR1A::::7.:C;MARK2::::7.:C;GRK4::::6.96:C;PDPK1::::6.96:C;PGFRB:::ant:6.96:DC;M4K3::::6.92:C;TNKS2::::6.92:C;ACK1::::6.92:C;KKCC1::::6.89:C;M3K7::::6.89:C;RET:M918T:::6.89:C;KCC2G::::6.85:C;M3K2::::6.85:C;CSF1R::::6.85:C;KIT:V559D-T670I::ant:6.82:DC;IKKE::::6.8:C;SIK1::::6.8:C;AURKC::::6.77:C;MARK1::::6.77:C;MINK1::::6.77:C;AAPK1::::6.74:C;IRAK3::::6.74:C;PGFRA:::ant:6.74:DC;PAK3::::6.74:C;LRRK2:G2019S:::6.74:C;PHKG1::::6.72:C;MAST1::::6.72:C;STK33::::6.72:C;KIT:V559D::ant:6.7:DC;M3K3::::6.68:C;KCC2B::::6.68:C;BMP2K::::6.66:C;KIT:::ant:6.66:DC;MYLK::::6.66:C;SLK::::6.66:C;HUNK::::6.62:C;KAPCB::::6.62:C;KS6A2::::6.62:C;KS6A5::::6.62:C;CSK21::::6.6:C;KGP1::::6.6:C;TYK2::::6.6:C;VGFR2:::ant:6.6:DC;KS6A1::::6.59:C;KS6A4::::6.59:C;ALK::::6.57:C;PI42B::::6.57:C;LCK::::6.55:C;MELK::::6.55:C;STK16::::6.55:C;KPCL::::6.54:C;PI51A::::6.51:C;NTRK2::::6.51:C;KPCD::::6.49:C;DYR1B::::6.48:C;SRPK2::::6.48:C;CLK1::::6.46:C;STK11::::6.46:C;RET::::6.46:C;TTK::::6.46:C;MARK4::::6.43:C;GAK::::6.42:C;NTRK1::::6.42:C;CLK4::::6.39:C;RIOK3::::6.38:C;ROS1::::6.37:C;VGFR1::::6.35:C;AAPK2::::6.34:C;BLK::::6.3:C;KPCE::::6.27:C;PIM1::::6.25:C;PIM3::::6.25:C;SIK2::::6.25:C;MET:Y1235D:::6.25:C;P3C2G::::6.24:C;LRRK2::::6.24:C;STK10::::6.23:C;UFO::::6.21:C;EGFR::::6.21:C;BRSK2::::6.19:C;M4K4::::6.19:C;MYLK4::::6.19:C;FAK2::::6.18:C;VGFR3::::6.17:C;JAK1::::6.17:C;KCC1D::::6.17:C;MET::::6.16:C;FGR::::6.14:C;HCK::::6.14:C;KPCA:::ant:6.14:DC;KAPCA::::6.14:C;KS6A3::::6.13:C;EGFR:L858R:::6.12:C;AKT2::::6.11:C;M3K10::::6.1:C;ABL1:T315I:::6.1:C;CLK2::::6.07:C;DAPK2::::6.05:C;PHKG2::::6.05:C;KPCT::::6.04:C;AKT1::::6.02:C;HIPK4::::6.02:C;MKNK2::::6.02:C;PRKX::::6.02:C;YES::::6.02:C;CDPK1::PLAF7::6.02:C;LATS1::::5.96:C;M4K5::::5.96:C;PK3CA:H1047L:::5.96:C;BRSK1::::5.92:C;FER::::5.92:C;RIOK1::::5.92:C;SRC::::5.92:C;CHK1::::5.89:C;ULK3::::5.89:C;KS6B1::::5.89:C;P3C2B::::5.85:C;TIE1::::5.85:C;SGK3::::5.85:C;KS6A6::::5.82:C;EGFR:G719C:::5.82:C;FGFR1::::5.8:C;TNIK::::5.8:C;KIT:V559D-V654A::ant:5.8:DC;FGFR3::::5.77:C;NTRK3::::5.77:C;DAPK3::::5.74:C;GSK3B::::5.74:C;STK25::::5.74:C;KCC1G::::5.74:C;ST17A::::5.72:C;TIE2::::5.72:C;KCC1A::::5.7:C;PAK1::::5.7:C;FYN::::5.68:C;M4K1::::5.68:C;PAK2::::5.68:C;MET:M1250T:::5.68:C;LATS2::::5.66:C;ERN1::::5.64:C;HIPK3::::5.64:C;ROCK2::::5.64:C;MYLK3::::5.64:C;FGFR2::::5.62:C;FRK::::5.62:C;ST32A::::5.62:C;GSK3A::::5.6:C;M4K2::::5.6:C;ZAP70::::5.59:C;M3K13::::5.55:C;EGFR:L861Q:::5.55:C;MERTK::::5.54:C;LTK::::5.52:C;EPHB6::::5.51:C;ERBB4::::5.51:C;HIPK2::::5.51:C;TBA1A::RAT::5.51:C;ABL1:H396P:::5.51:C;PIM2::::5.51:C;KPCD3::::5.49:C;MK10::::5.44:C;CLK3::::5.44:C;DMPK::::5.42:C;IKKA::::5.42:C;LYN::::5.38:C;MK08::::5.36:C;AKT3::::5.36:C;WEE1::::5.34:C;DAPK1::::5.33:C;ST17B::::5.33:C;DUSTY::::5.33:C;MP2K4::::5.32:C;TSSK1::::5.32:C;MK09::::5.3:C;MP2K3::::5.28:C;EGFR:G719S:::5.28:C;ICK::::5.23:C;KPCD2::::5.2:C;IKKB::::5.2:C;MP2K6::::5.19:C;E2AK2::::5.16:C;CDK19::::5.14:C;DDR1::::5.14:C;ROCK1::::5.11:C;CSK::::5.06:C|CP343:::ind::D;CP3A7:::ind::D;CP3A5:::ind::D;CP3A4:::duo::D;CP2E1:::inh::D;CP2D6:::inh::D;CP2CJ:::duo::D;CP2C9:::duo::D;CP2C8:::duo::D;CP2B6:::ind::D;CP1A2:::duo::D;CP3A4,CP343,CP3A5,CP3A7:::duo::D||
Nemonoxacin|inv||CP1A2:::inh::D||
Reslizumab|ok_inv|IL5:::ant::D|||
Panobinostat|ok_inv|HDAC4::::9.22:C;HDAC2::::9.19:C;HDAC5::::9.15:C;HDAC6::::9.15:C;HDAC1,HDA10,HDA11,HDAC2,HDAC3,HDAC4,HDAC5,HDAC6,HDAC7,HDAC8,HDAC9:::inh:9.08,8.4,8.46,9.19,8.96,9.22,9.15,9.15,8.64,8.31,8.92:DC;HDAC1::::9.08:C;HDAC3::::8.96:C;HDAC9::::8.92:C;HDAC7::::8.64:C;HDA11::::8.46:C;HDA10::::8.4:C;HDAC8::::8.31:C|CP3A4:::sub::D;CP2D6:::inh::D|MDR1:::sub::D|
Apixaban|ok|FA10:::inh:10.1:DC;FA10::RABIT::9.77:C;THRB::::5.51:C|CP3A5:::sub::D;CP2J2:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP1A2:::sub::D;CP3A4:::sub::D|ABCG2:::sub::D;MDR1:::sub::D|
Catumaxomab|ok_out|EPCAM:::lig::D;FCG2A:::ago::D;FCG3A:::ago::D;FCG3B:::ago::D;CD3E:::ago::D;FCGR1:::ago::D|||
Tafenoquine|ok_inv||FENR::PLAF7:sub::D;CP2D6:::sub::D|S47A2:::inh::D;S47A1:::inh::D;S22A2:::inh::D|
Mepolizumab|ok_inv|IL5:::ant::D|||
Peramivir|ok_inv|NRAM::I18A0::9.08:C;NRAM::I34A1::8.85:C;NRAM::INBLE::8.3:C;NRAM::INBBE:::D;NRAM::I79A0:::D;NRAM::I75A5:::D|||
Bosutinib|ok|ABL1:F317L::inh:10.54:DC;ABL1:Y253F::inh:10.44:DC;ABL1:M351T::inh:10.43:DC;ABL1:Q252H::inh:10.41:DC;ABL1:E255K::inh:10.33:DC;ABL1:H396P::inh:10.24:DC;ABL1:::inh:10.24:DC;ABL1:F317I::inh:9.74:DC;M4K5::::9.52:C;YES::::9.4:C;ABL2::::9.3:C;LCK::::9.23:C;ERBB3::::9.11:C;MP2K1:::inh:9.:DC;SRC:::inh:9.:DC;BMX::::9.:C;FGR::::8.96:C;GAK::::8.89:C;FRK::::8.85:C;FYN::::8.74:C;STK35::::8.7:C;BTK::::8.6:C;ACK1::::8.57:C;M4K2::::8.51:C;MINK1::::8.49:C;HCK:::inh:8.49:DC;BLK::::8.48:C;ABL1:T315I::inh:8.44:DC;STK24::::8.41:C;LYN::::8.38:DC;SLK::::8.33:C;M4K3::::8.29:C;EPHB4::::8.26:C;EPHA3::::8.24:C;STK10::::8.15:C;BLK::MOUSE::8.14:C;MP2K5::::8.09:C;M4K4::::8.09:C;EPHB2::::8.08:C;EPHA8::::8.05:C;MP2K2:::inh:8.:DC;M4K1::::7.82:C;M3K19::::7.8:C;EGFR::::7.74:C;EPHA2::::7.74:C;EPHA4::::7.74:C;NTRK1::::7.66:C;EGFR:L858R:::7.64:C;EGFR:G719S:::7.59:C;ERBB4::::7.59:C;EPHA5::::7.57:C;NTRK2::::7.57:C;SIK2::::7.54:C;M3K2:::inh:7.52:DC;SIK1::::7.52:C;TNIK::::7.51:C;CSK::::7.49:C;EPHB1::::7.48:C;STK26::::7.43:C;STK33::::7.43:C;TXK::::7.4:C;IKKE::::7.28:C;UFO::::7.28:C;KSYK::::7.28:C;M3K3::::7.27:C;TYRO3::::7.21:C;SIK3::::7.19:C;EGFR:L861Q:::7.15:C;KIT:D816V:::7.14:C;M3K20::::7.1:C;DMPK::::7.04:C;KCC1D::::7.04:C;WEE2::::7.03:C;EGFR:G719C:::7.01:C;SRMS::::7.:C;M3K7::::7.:C;M3K4::::6.96:C;MERTK::::6.96:C;KC1E::::6.96:C;CHK2::::6.92:C;DDR1::::6.92:C;HIPK4::::6.89:C;KIT:V559D-V654A:::6.89:C;FAK2::::6.87:C;DDR2::::6.85:C;ALK:L256T:::6.82:C;TNI3K::::6.77:C;KIT:D816H:::6.74:C;KCC2G:::inh:6.74:DC;STK4::::6.72:C;PGFRB::::6.7:C;EPHB3::::6.68:C;NUAK2::::6.66:C;KC1D::::6.62:C;TBK1::::6.6:C;E2AK4::::6.57:C;KIT:A829P:::6.57:C;KC1A::::6.55:C;TEC::::6.55:C;CLK3::::6.52:C;FES::::6.48:C;EGFR:T790M:::6.47:C;PHKG1::::6.47:C;TAOK3::::6.47:C;MAST1::::6.46:C;BMP2K::::6.46:C;PMYT1::::6.46:C;FER::::6.44:C;IRAK4::::6.44:C;ROCK2::::6.44:C;STK3::::6.43:C;DUSTY::::6.42:C;CSF1R::::6.42:C;EGFR:L858R-T790M:::6.41:C;KIT::::6.38:C;KIT:V559D:::6.37:C;ULK2::::6.35:C;ULK3::::6.34:C;M3K13::::6.32:C;MYLK::::6.31:C;ERBB2:T790M:::6.31:C;LRRK2::::6.3:C;WEE1::::6.29:C;HIPK1::::6.28:C;KIT:L576P:::6.28:C;FAK1::::6.27:C;TLK1::::6.24:C;STK36::::6.24:C;BMPR2::::6.24:C;IRAK1::::6.22:C;CLK1::::6.22:C;E2AK1::::6.2:C;NEK11::::6.19:C;KS6B1::::6.18:C;M3K12::::6.17:C;ALK::::6.16:C;VRK2::::6.15:C;KKCC2::::6.11:C;LRRK2:G2019S:::6.08:C;CSKP::::6.08:C;ROCK1::::6.06:C;STK25::::6.05:C;KPCT::::6.04:C;PLK2::::6.02:C;FLT3:D835H:::6.:C;EPHA6::::5.96:C;FLT3:D835Y:::5.96:C;JAK2::::5.96:C;JAK3::::5.92:C;CDK7::::5.92:C;ULK1::::5.92:C;KS6A3::::5.92:C;TIE2::::5.92:C;TAOK1::::5.89:C;PHKG2::::5.89:C;MP2K6::::5.89:C;CDK14::::5.85:C;NIM1::::5.82:C;KPCD::::5.8:C;CDK15::::5.8:C;ZAP70::::5.8:C;NEK2::::5.8:C;RIOK3::::5.8:C;ITK::::5.77:C;GRK7::::5.77:C;CLK2::::5.77:C;ST32A::::5.74:C;PLK1::::5.74:C;TAOK2::::5.72:C;HIPK2::::5.72:C;PAK2::::5.72:C;ANKK1::::5.68:C;TLK2::::5.68:C;NLK::::5.66:C;RIOK1::::5.66:C;MET::::5.66:C;FLT3::::5.66:C;FLT3:K663Q:::5.66:C;EPHA1::::5.64:C;AAK1::::5.64:C;MYO3B::::5.64:C;PAK1::::5.64:C;MK07::::5.64:C;CTRO::::5.62:C;KPCE::::5.62:C;CDK16::::5.62:C;ERBB2::::5.6:C;KC1AL::::5.59:C;MP2K3::::5.59:C;MP2K4::::5.59:C;KS6A6::::5.57:C;M3K9::::5.57:C;M3K11::::5.57:C;TIE1::::5.54:C;PKN1::::5.54:C;CHK1::::5.52:C;EPHB6::::5.52:C;LTK::::5.52:C;MET:Y1235D:::5.51:C;HIPK3::::5.49:C;PKN2::::5.49:C;KS6A2::::5.49:C;CLK4::::5.49:C;PI51A::::5.48:C;NTRK3::::5.47:C;FLT3:N841I:::5.47:C;STK39::::5.43:C;RIPK2::::5.43:C;RET:M918T:::5.42:C;SRPK3::::5.41:C;AAPK1::::5.41:C;PGFRA::RAT::5.4:C;RET:V804M:::5.38:C;M3K1::::5.36:C;KCC2A::::5.35:C;TYK2::::5.35:C;KPCD3::::5.34:C;TSSK1::::5.34:C;RET::::5.32:C;GRK4::::5.31:C;HUNK::::5.3:C;PGFRA::::5.29:C;MP2K7::::5.28:C;DCLK3::::5.27:C;PKNB::MYCTU::5.26:C;MATK::::5.24:C;PAK3::::5.24:C;NUAK1::::5.23:C;MYO3A::::5.21:C;RON::::5.2:C;MET:M1250T:::5.17:C;CDK2:::inh::D;BCR:::inh::D|CP2C8:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Flupirtine|inv|NFKB1::::7.55:C;HIF1A::::5.4:C;CP3A4::::5.1:C;CASP7::::5.:C;ADA2A|||
Axitinib|ok_inv|VGFR2:::inh:9.6:DC;ABL1::::9.38:C;KIT:V559D:::9.31:C;PGFRA::::9.29:C;PGFRB::::9.24:C;AURKC::::8.89:C;KIT:V559D-T670I:::8.85:C;ABL1:T315I:::8.82:C;KIT:L576P:::8.77:C;KIT::::8.49:C;KIT:V559D-V654A:::8.46:C;VGFR2:E990V::inh:8.42:DC;PLK4::::8.38:C;VGFR1:::inh:8.24:DC;AURKB::::7.96:C;ABL1:H396P:::7.7:C;CSF1R::::7.68:C;FLT3:K663Q:::7.51:C;ABL1:M351T:::7.44:C;FLT3::::7.38:C;FGFR1::::7.25:C;ABL1:E255K:::7.2:C;ABL2::::7.15:C;AURKA::::7.14:C;TIE1::::7.01:C;RET:M918T:::7.:C;FGFR2::::6.96:C;RET::::6.92:C;MP2K5::::6.85:C;TNK1::::6.8:C;VGFR3:::inh:6.77:DC;TNIK::::6.74:C;ABL1:Q252H:::6.7:C;FLT3:N841I:::6.7:C;FGFR3::::6.68:C;FGFR3:G697C:::6.68:C;ABL1:Y253F:::6.64:C;M3K19::::6.57:C;FLT3:D835Y:::6.57:C;TIE2::::6.51:C;ABL1:F317L:::6.48:C;M4K1::::6.48:C;FLT3:D835H:::6.48:C;DDR1::::6.47:C;M4K4::::6.46:C;EPHB6::::6.44:C;STK16::::6.43:C;UFO::::6.38:C;CDKL2::::6.28:C;M4K5::::6.26:C;MINK1::::6.25:C;ULK3::::6.17:C;ABL1:F317I:::6.1:C;MET::::6.09:C;LRRK2::::6.04:C;SLK::::6.:C;BMP2K::::6.:C;LRRK2:G2019S:::6.:C;MET:Y1235D:::6.:C;RIOK3::::6.:C;MET:M1250T:::5.96:C;MK10::::5.96:C;CSK::::5.96:C;ITK::::5.92:C;STK10::::5.92:C;AAK1::::5.92:C;RIOK1::::5.92:C;M4K3::::5.92:C;M4K2::::5.89:C;RET:V804L:::5.89:C;NUAK2::::5.89:C;MYLK2::::5.89:C;KIT:D816V:::5.89:C;STK4::::5.85:C;RIPK4::::5.85:C;KKCC1::::5.85:C;KKCC2::::5.82:C;HUNK::::5.82:C;RET:V804M:::5.8:C;M3K12::::5.77:C;MYLK3::::5.77:C;FGR::::5.74:C;KIT:A829P:::5.74:C;NTRK1::::5.74:C;SRPK1::::5.74:C;MYO3A::::5.72:C;SIK1::::5.68:C;STK3::::5.66:C;EGFR:G719C:::5.64:C;SRPK3::::5.64:C;GRK4::::5.64:C;TXK::::5.62:C;FLT3:R834Q:::5.62:C;RIPK1::::5.6:C;MP2K2::::5.59:C;M3K20::::5.59:C;GAK::::5.57:C;LCK::::5.57:C;YES::::5.57:C;PKN2::::5.57:C;MP2K1::::5.57:C;CSK22::::5.55:C;M3K3::::5.55:C;BMR1B::::5.54:C;M3K9::::5.52:C;JAK3::::5.51:C;IRAK1::::5.51:C;BLK::::5.51:C;MERTK::::5.49:C;ROS1::::5.49:C;JAK2::::5.48:C;ANKK1::::5.44:C;TYK2::::5.44:C;MK08::::5.41:C;TTK::::5.41:C;KIT:D816H:::5.38:C;TESK1::::5.37:C;PAK4::::5.35:C;MRCKB::::5.32:C;CDK16::::5.28:C;DDR2::::5.28:C;AVR2B::::5.28:C;M3K4::::5.25:C;ACK1::::5.22:C;EGFR:G719S:::5.21:C;E2AK2::::5.13:C;ULK2::::5.:C;RIPK2::::5.:C|UD11:::sub::D;CP2CJ:::sub::D;CP1A2:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|SO1B1:::inh::D;MDR1:::sub::D|
Casopitant|inv|NK1R::::9.9:DC;SGMR1::::5.53:C;CP3A4::::5.31:DC|||
Isavuconazonium|ok_inv||CP3A4:::duo::D|MDR1:::inh::D|
Dalfampridine|ok|CP2D6::::7.2:C;TSHR::::6.9:C;LMNA::::6.05:C;CYSP::TRYCR::5.5:C;LEF::BACAN::5.1:C;TAU::::5.05:C;MK01::::5.:C;KCND3:::ant::D;KCND2:::ant::D;KCND1:::ant::D;KCNC3:::ant::D;KCNC2:::ant::D;KCNC1:::ant::D;KCNB2:::ant::D;KCNB1:::ant::D;KCA10:::ant::D;KCNA7:::ant::D;KCNA6:::ant::D;KCNA5:::ant::D;KCNA4:::ant::D;KCNA3:::ant::D;KCNA2:::ant::D;KCNA1:::ant::D|CP2E1:::sub::D|S22A2:::sub::D|
Denosumab|ok|TNF11:::abo::D|||
Ofatumumab|ok|CD20:::inh::D|||
Safinamide|ok_inv|AOFB:::ant:8.29:DC;AOFB::RAT::7.74:C|CP3A5:::inh::D;CP2E1:::inh::D;CP2CJ:::inh::D;CP2D6:::inh::D;CP2C9:::inh::D;CP2B6:::inh::D;CP1A2:::inh::D;CP1A1:::inh::D;CP3A4:::sub::D;AOFA:::inh::D|SO3A1:::sub::D;ABCG2:::inh::D|
Liraglutide|ok|GLP1R:::ago::D|DPP4:::sub::D;NEP:::sub::D||ALBU:::bin::D
Abetimus|inv||||
Pasireotide|ok|SSR1;SSR2;SSR3;SSR5|CP3A4:::inh::D||
Golimumab|ok|TNFA:::abo::D|||
Belatacept|ok_inv|CD86:::ant::D;CD80:::ant::D|||
Naproxcinod|inv||||
Clevudine|inv||||
Vilazodone|ok|5HT1A:::ago:9.52:DC;5HT1A::RAT::9.52:C;SC6A4::RAT::9.3:C;SC6A4:::inh:9.3:DC;DRD3::RAT::7.15:C;5HT4R::RAT::6.6:C;DRD2::RAT::6.18:C;DRD2::::6.18:C;5HT2A::RAT::5.82:C;5HT2C::RAT::5.7:C;ADA1A::::5.7:C;5HT6R::RAT::5.52:C;5HT7R::RAT::5.52:C;DRD4::RAT::5.47:C;5HT1D::RAT::5.4:C;5HT3A::RAT::5.37:C;5HT1B::RAT::5.3:C;ADA2A::::5.22:C|CP2CJ:::sub::D;CP2D6:::sub::D;CP3A4:::sub::D||
Laquinimod|inv||CP3A4:::sub::D||
Sipuleucel_T|ok_inv|PPAP|||
Ethanolamine_oleate|ok|Calcium_ions:::chel::D;FA12:::act::D|||
Nitrous_oxide|ok_vet||||
Mepyramine|ok_vet|HRH1:::ant:10.85:DC;HRH1::CAVPO::9.5:C;LMNA::::8.96:C;AA3R::::8.89:C;HRH1::RAT::8.24:C;SC6A4::::7.6:C;5HT2A::::6.55:C;5HT2C::::6.23:C;CP3A4::::6.2:C;SGMR1::::6.18:C;SC6A3::::6.16:C;KCNH2::::5.96:C;ADA2A::::5.95:C;5HT2B::::5.75:C;TSHR::::5.3:C;CP2CJ::::5.:C|CP2D6:::inh:7.:DC|S22A5;S22A4|
Aprotinin|ok_out|TRY1;CTRB1;PLMN;KLK1|CHLE:::inh::D||
Xylometazoline|ok_inv|5HT1D::::9.15:C;ADA1B::RAT::8.32:C;5HT1B::::7.89:C;ADA2C::RAT::7.64:C;ADA1A:::ago:7.04:DC;P53::::5.5:C;TSHR::::5.4:C;CP2D6::::5.4:C;ACM1::RAT::5.25:C;LMNA::::5.1:C;ADA2C:::ago::D;ADA1D:::ago::D;ADA1B:::ago::D;ADA2B:::ago::D;ADA2A:::ago::D|||
Dabigatran_etexilate|ok|THRB:::inh:8.58:DC|NQO2:::inh::D;UDB15:::sub::D;UD2B7:::sub::D;UD19:::sub::D;EST2:::sub::D;EST1:::sub::D|MDR1:::sub::D|
Arbekacin|exp_inv|RS12::ECOLI:inh::D|||
Artemether|ok|LMNA::::6.25:C|CP2CJ:::sub_ind::D;CP2C9:::sub::D;CP2B6:::sub_ind::D;CP3A5:::sub::D;CP3A4:::sub_ind::D||
Betahistine|ok_inv|HRH3::RAT::5.69:C;HRH3:::ant::D;HRH1:::ago::D|||
Degarelix|ok|GNRHR:::ant:9.24:DC|||
Desvenlafaxine|ok_inv|SC6A4:::inh:7.82:DC;ADA1A::RAT::7.22:C;SC6A4::RAT::6.74:C;SC6A2:::inh:5.82:DC;SC6A3:::inh::D|CP2D6:::inh::D;CP3A4:::inh::D||
Dexmethylphenidate|ok_inv|SC6A3:::inh:7.8:DC;SC6A3::RAT::7.62:C;SC6A4:::inh::D;SC6A2:::inh::D|Carboxylesterase::ALCSP:sub::D||
Fesoterodine|ok|ACM5:::ant::D;ACM2:::ant::D;ACM1:::ant::D;ACM4:::ant::D;ACM3:::ant::D|CP2D6:::sub::D;CP3A4:::sub::D|MDR1:::sub::D|
Gadobutrol|ok||||
Iobenguane|ok_inv|TPO::::5.8:C||SC6A2:::sub::D|
Gadofosveset_trisodium|ok||||ALBU:::sub::D
Isometheptene|ok|ADA1A:::ago::D;VMAT2:::inh::D|||
Levonordefrin|ok|ADA2C::RAT::8.11:C;HCD2::::7.:C;LMNA::::6.6:C;TYDP1::::6.45:C;HIF1A::::6.3:C;ADA1B::RAT::6.11:C;RECQ1::::5.75:C;KPYK::LEIME::5.5:C;LOX15::::5.5:C;KDM4E::::5.35:C;ADA2A,ADA2B,ADA2C:::ago::D|||
Lumefantrine|ok||CP2D6:::inh::D;CP3A4:::sub_ind::D||
Methacholine|ok_inv|ACM2::RAT::7.23:C;ACM2::::7.23:C;ACM3::RAT::6.92:C;ACM1::RAT::6.4:C;ACM4::RAT::6.15:C;ACM4::::5.8:C;ACM3:::ago::D|||
Methyltestosterone|ok|ANDR::RAT::8.37:C;GCR::::6.08:C;ESR1;ANDR:::ago::D|CP19A:::sub_ind::D;CP3A4:::sub::D;CP2B6:::sub::D|S22A8:::ind::D;SO1A2:::duo::D|SHBG::::8.43:DC;ALBU
Naphazoline|ok_inv|ADA2C::::8.64:C;ADA2C::RAT::8.32:C;ADA1B::RAT::8.24:C;ADA1A:::ago:7.2:DC;NISCH::::6.92:C;NISCH::RAT::6.61:C;TAU::::6.1:C;LMNA::::5.7:C;MK01::::5.4:C;CP2D6::::5.1:C;ADA2A:::ago::D|||
Nilvadipine|ok_inv|CAC1C::RAT::8.98:C;NR1I2::::6.05:C;CA2D3:::inh::D;CAC1S:::inh::D;CAC1D:::inh::D;CACB2:::inh::D;CA2D1:::inh::D;CAC1C:::inh::D|CP2E1:::sub::D;CP2C8:::inh::D;CP2CJ:::inh::D;CP2A6:::inh::D;CP3A4:::inh::D||
Norelgestromin|ok_inv|ANDR:::pag::D;ALBU;PRGR:::ago::D|CP3A4:::sub::D;STS:::inh::D||
Propylhexedrine|ok|VMAT2;TAAR1:::ago::D|||
Potassium_Iodide|ok|Tyrosine:::bin::D|||
Fospropofol|ok_ill_inv|GBRB2:::pot::D;GBRB3:::pot::D|PPBT:::sub::D||ALBU:::sub::D
Fosaprepitant|ok||CP3A4:::duo::D;CP2C9:::ind::D||
Stanozolol|ok_vet|ANDR::RAT::7.82:C;ESR1::::7.49:C;CP2CJ::::7.32:C;CP2C9::::5.95:C;AA3R::::5.33:C;CP2D6::::5.03:C;Glucocorticoid_binding_proteins:::bin::D;ANDR:::ago::D|||
Buserelin|ok_inv|LSHR;GNRHR|CP19A:::ind::D||
Velaglucerase_alfa|ok_inv|GLCM|||
Aluminum_hydroxide|ok_inv||||
Calcium_carbonate|ok_inv||||
Lornoxicam|ok_inv|AMPC::ECOLI::5.1:C;PGH2:::inh::D;PGH1:::inh::D|CP2C9:::sub::D||
Sparteine|exp||CP2D6:::inh::D||
Sulfaphenazole|ok|ACM1::RAT::7.65:C;CP3A4::::6.9:C;DPOLB::::6.05:C;NPSR1::::5.5:C;TSHR::::5.4:C;NFKB1::::5.15:C;LMNA::::5.1:C;HCD2::::5.:C;DHPS::ECOLI:inh::D|CP2C9:::inh:7.3:DC;CP2D6:::inh::D;CP2C8:::inh::D;CP2B6:::inh::D||
Gestodene|inv|PRGR:::bin::D|CP2CJ:::inh::D;CP3A4:::sub::D;CP3A7:::inh::D;CP3A5:::inh::D||
Aceclofenac|ok_inv|LMNA::::7.35:C;TTHY::::5.92:C;ALDR::RAT::5.89:C;UBP2::::5.5:C;KMT2A::::5.45:C;MK01::::5.23:C;PGH1:::inh::D;PGH2:::inh::D|CP2C9:::sub:5.8:DC||
Ketobemidone|inv|SGMR1::RAT::8.7:C;OPRM::MOUSE::5.15:C;NMDA:::ant::D;OPRD:::ago::D;OPRK:::ago::D;OPRM:::ago::D|CP2C8:::sub::D;CP2CJ:::sub::D;CP2B6:::sub::D;UD19:::sub::D;CP3A4:::sub::D;CP2C9:::sub::D;PGH1:::sub::D||
Seratrodast|exp|TA2R:::ant:8.13:DC|CP2A6:::inh::D;PGH1:::sub::D;UD19:::sub::D;CP2B6:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP3A4:::sub_ind::D;CP2C9:::sub::D||
Ambroxol|ok_inv|CP2D6::::6.25:C;SC6A4::::5.74:C;GLCM::::5.39:C|CP3A4:::sub::D||
Drotaverine|ok_inv|PDE4A:::inh::D;CAC1C:::inh::D|||
Chymopapain|ok_out|PRG2:::degr::D|||
Triclofos|ok_out||||
Danaparoid|ok_out|ANT3:::aga::D|||
Beta_carotene|ok_nutra|SO1B1::::6.47:C;SO1B3::::5.65:C;Free_radicals:::bin::D|BCDO1:::sub::D||RET5:::sub::D;RET4:::sub::D;RET3:::sub::D;RET2:::sub::D;RET1:::sub::D;VLDLR:::sub::D
Glycine_betaine|ok_nutra|TSHR::::8.4:C;BCL2|PROD:::inh::D;CHLE:::inh::D||
Manganese|ok_nutra|IDH3A;IDH3G;TAB1;ARGI1;TRFE|ACOC:::inh::D||
Fomivirsen|ok_out|VIE3::HCMVT:oli::D;IE247::HCMVT:oli::D|||
Sacrosidase|ok||||
Beractant|ok||||
Pinacidil|ok|KCJ11::::6.49:C;AMPC::ECOLI::6.45:C;LMNA::::5.9:C;AGAL::::5.5:C;BLM::::5.45:C;ABCC9::::5.45:C;NPSR1::::5.3:C|CP3A4:::sub:5.5:DC||
Tetryzoline|ok|ADA1B::RAT::7.96:C;ADA2C::RAT::7.52:C;ADA1A:::ago::D|||
Alcaftadine|ok|HRH1:::ant::D|||
Ammonium_chloride|ok_inv_vet||||
Ammonium_lactate|ok||||
Bendamustine|ok_inv|HDAC6::::8.22:C;HDAC2::::8.05:C;HDAC1::::7.77:C;HDAC3::::7.6:C;HDA10::::7.14:C;HDAC8::::6.97:C|CP1A2:::sub::D||
Benzyl_alcohol|ok|TSHR::::7.7:C|CP2D6:::sub::D;CP2E1:::sub::D;CP1A2:::sub::D;ALDH2:::sub::D;CP1A1:::inh::D;CP2C8:::sub::D||
Besifloxacin|ok|PARC::HAEIN:ant::D;PARC::STRPN:ant::D;GYRA::HAEIN:ant::D;GYRA::STRPN:ant::D|CP1A2:::inh::D||
Cabazitaxel|ok|TBA4A:::bin::D;TBB1:::bin::D|CP3A4:::sub::D;CP3A5:::sub::D;CP2C8:::sub::D|MDR1:::inh::D;ABCG2:::inh::D;SO1B1:::inh::D;SO1B3:::inh::D|
Human_calcitonin|ok_inv|ACTN1:::destbz::D|ANAG:::sub::D;AMPN:::sub::D;PGM1:::sub::D||
Capsaicin|ok|TRPV1:::ago:8.6:DC;TRPV1::RAT::7.72:C;TRPV4::RAT::7.52:C;PGH1::::5.81:C;AL1A1::::5.7:C;PHB2|CP3A4:::inh:5.6:DC;CP1A2:::sub_ind:5.52:DC;CHLE:::inh::D;GLNA:::ind::D;DOPO:::inh::D;AOFA:::inh::D;CP2E1:::sub::D;PERM:::inh::D;PGH2:::inh::D||
Carglumic_acid|ok|CPSM:::alo::D|||
Sodium_cellulose_phosphate|ok|Calcium_ions:::bin::D|||
Chenodeoxycholic_acid|ok|NTCP2::::5.48:C;NR1H4::::5.47:DC;GPBAR::::5.21:DC;AK1C2:::sub::D;NR1I2|UD2B7:::inh::D;CP3A4:::sub::D;CP27A:::sub::D||
Cupric_sulfate|ok||PH4H:::ind::D;LYOX:::ind::D;COX1:::ind::D|ALBU;CERU|
Dalteparin|ok|ANT3:::pot::D;VEGFA:::inh::D;TFPI1:::inh::D;LYAM3:::inh::D|HPSE:::sub::D||
Desoxycorticosterone_acetate|ok|TAU::::6.75:C;LMNA::::5.4:C;MCR:::ago::D|CP3A4:::sub::D||
Difluprednate|ok|HIF1A::::8.4:C;LMNA::::6.25:C;NPSR1::::5.6:C;GCR:::ago::D|CP3A4:::sub::D||
Dimercaprol|ok|AL1A1::::7.:C;HCD2::::6.:C;FFP::BACIU::5.65:C;CP1A2::::5.4:C;NR1I2::::5.3:C;A4;Mercury:::chel::D;Cadmium:::chel::D;Arsenic:::chel::D|||
Prussian_blue|ok||||
Gallium_citrate_Ga_67|ok|||TFR1:::sub::D;Q19KS1:::sub::D;FRIL:::sub::D;FRIH:::sub::D|
Ganirelix|ok|GNRHR:::ant:9.3:DC|||
Halcinonide|ok_out|GCR::::9.14:C;ANDR::RAT::6.23:C;AMPC::ECOLI::5.:C;SMO:::ago::D|CP3A4:::sub::D||
Hexocyclium|ok|ACM1:::ant::D;ACM2:::ant::D;ACM3:::ant::D;ACM4:::ant::D|||
Histrelin|ok|GNRHR:::ago::D|||
Hydroxyprogesterone_caproate|ok_inv|DNAB::MYCTU::5.69:C;HIF1A::::5.4:C;RECA::MYCTU::5.31:C;NPSR1::::5.:C;HD::::5.:C;PRGR:::ago::D|CP2CJ:::ind::D;CP3A5:::sub::D;CP3A4:::sub::D||
Lanreotide|ok|SSR2:::ago:9.3:DC;SSR5:::ago:8.4:DC;SSR3::::7.2:C;SSR1::::6.3:C|CP3A4:::inh::D||
Lanthanum_carbonate|ok|Phosphate:::bin::D|||
Lodoxamide|ok||||
Mafenide|ok_vet|CAH12::::9.52:C;CAH13::MOUSE::7.39:C;CAH7::::7.12:C;CAH9::::6.99:C;CAH2::::6.77:C;CAN::CANAL::6.77:C;CAH::METTE::6.46:C;CAN::YEAST::6.36:C;CYNT::HELPY::6.08:C;CAH15::MOUSE::6.01:C;CAH4::BOVIN::5.55:C;CAH4::::5.55:C;CAH14::::5.49:C;CAH6:::ant:5.32:DC;MTCA1::MYCTU::5.06:C|||
Mangafodipir|ok_out||SODM:::act::D|NRAM2:::sub::D|A2MG:::bin::D;ALBU:::bin::D
Mebutamate|ok||||
Methenamine|ok_vet||||
Methylnaltrexone|ok|OPRM:::ant::D;OPRK:::ant::D|||
Nepafenac|ok_inv|PGH2:::inh::D;PGH1:::inh::D|||
Niclosamide|ok_inv_vet|ACM1::RAT::8.74:C;LMNA::::7.6:C;NPC1::::7.4:C;RAB9A::::7.1:C;TPO::::7.:C;SMN::::6.9:C;LEF::BACAN::6.6:C;STAT3::::6.6:C;GEMI::::6.5:C;PMP22::::6.42:C;CP2CJ::::6.4:C;P53::::6.3:C;TSHR::::6.3:C;RORG::MOUSE::6.25:C;LUCI::PHOPY::6.1:C;HD::::6.1:C;MTOR::::5.93:C;HIF1A::::5.7:C;CP3A4::::5.6:C;KPYK::LEIME::5.6:C;MEN1::::5.55:C;TAU::::5.5:C;KPYM::::5.5:C;AL1A1::::5.45:C;CYSP::TRYCR::5.25:C;AMPC::ECOLI::5.25:C;SRC::::5.:C;JAK2::::5.:C;DNA:::ant::D|CP2C9:::sub:6.2:DC;CP1A2:::inh:5.9:DC||
Nonoxynol_9|ok_out|LMNA::::8.05:C;SO1B1::::5.72:C;SO1B3::::5.54:C;MEN1::::5.15:C;CYSP::TRYCR::5.:C|PGH2:::ind::D||
Phenyl_aminosalicylate|ok|LMNA::::6.05:C;TAU::::5.5:C;P53::::5.:C|||
Plerixafor|ok|CCR2::::10.4:C;CXCR4:::ant:9.09:DC;CXCR4::RAT::7.:C|||
Plicamycin|ok_out|DNA:::ant::D|||
Polidocanol|ok|THB::::7.05:C|||
Povidone_iodine|ok||||
Pralatrexate|ok_inv|TYSY:::inh::D;DYR:::inh::D|FOLC:::sub::D|S19A1:::sub::D|
Protokylol|ok_vet|ADRB2:::ago::D|||
Pyrithione|ok|RORG::MOUSE::7.2:C;LMNA::::7.:C;LOX15::::6.7:C;LEF::BACAN::6.4:C;HD::::6.05:C;CYSP::TRYCR::6.:C;AL1A1::::5.9:C;HCD2::::5.9:C;P53::::5.6:C;HIF1A::::5.5:C;TYDP1::::5.3:C;TSHR::::5.2:C;PGDH::::5.:C|||
Pyrvinium|ok||||
Raltegravir|ok|CCR1::::8.3:C;Integrase::9HIV1:inh::D|UD11:::sub::D||
Phenylbutyric_acid|ok_inv|HDAC1::::5.55:C;THER::BACTH:::D;TYRB::PARDE:::D|CP2D6:::inh::D||
Sulconazole|ok|CP2CJ::::7.8:C;CP3A4::::7.15:C;SC6A4::::7.12:C;THAS::::6.74:C;ACM4::::6.26:C;ACM3::::6.14:C;ADA2C::::6.14:C;ACM1::::6.05:C;DRD3::::5.98:C;5HT2A::::5.95:C;SC6A3::::5.86:C;5HT2C::::5.84:C;AA3R::::5.83:C;ADA2A::::5.82:C;ADA2B::::5.79:C;NK2R::::5.78:C;ACM5::::5.73:C;5HT2B::::5.72:C;SC6A2::::5.7:C;FYN::::5.43:C;I23O1::::5.19:C;NR1H4::::5.16:C;I23O2::MOUSE::5.:C|CP2C9:::inh:6.7:DC;CP1A2:::inh:6.22:DC;CP2D6:::inh:6.1:DC||
Sulfameter|ok|AMPC::ECOLI::6.45:C;DHPS::ECOLI:inh::D|||
Tinzaparin|ok|ANT3:::pot::D;ITA4:::inh::D;SDF1:::bin::D|ATS4:::inh::D||
Tiopronin|ok_inv|TYDP1::::6.:C;ACE::RABIT::5.72:C|PERM:::inh::D||
Triethylenetetramine|ok_inv|LMNA::::6.3:C||GPC1::BOVIN:sub::D|
Triptorelin|ok_vet|GNRHR:::ago::D|||
Unoprostone|ok_inv||||
Viomycin|ok|TLYA::MYCTU:inh::D|||
Hymecromone|exp_inv|LMNA::::8.35:C;CAH9::::6.25:C;DHB3::::6.:C;HCD2::::5.6:C;CP1A2::::5.4:C;CAH12::::5.09:C;Arylsulfate_sulfotransferase_AssT::ECOK1:::D|||
Azapropazone|out||||ALBU
Felbinac|exp|PGH1::::6.05:C;LMNA::::5.6:C;TSHR::::5.3:C;CATL1|||
Chloramphenicol_succinate|ok|DRAA::ECOLX:::D|||
Dibromotyrosine|exp|AL1A1::::5.4:C;HCD2::::5.2:C;EPOR|||
Flavone|ok_exp|P53::::8.3:C;CP19A::::8.1:C;GBRA1::::7.77:C;TNKS2::::6.85:C;TNKS1::::6.49:C;GBRP::RAT::6.:C;PARP1::::5.86:C;CAH1::::5.73:C;RAB9A::::5.5:C;AA1R::RAT::5.48:C;AA2AR::RAT::5.46:C;AA2BR::RAT::5.46:C;CAH9::::5.38:C;NPC1::::5.25:C;ANDR::::5.23:C;CAH12::::5.14:C;CAH2::::5.06:C;PGDH::::5.05:C;CP1B1;ERR2:::ago::D;ERR1:::ago::D;NCZS::STRCZ:::D|||
Fasudil|inv|ROCK1::::7.5:DC;ROCK2::::7.3:DC;PRKX::::7.3:C;KAPCA::::7.1:DC;CP2D6::::6.7:C;CLK4::::6.5:C;KAPCB::::6.34:C;KPCT::::6.2:C;PKN2::::6.11:C;KS6A3::::6.:C;KS6B1::::6.:C;KPCD3::::6.:C;CDK8::::5.9:C;KPCD2::::5.9:C;DAPK3::::5.9:C;PKN1::::5.77:C;ROCK2::RAT::5.72:C;LRRK2::::5.7:C;CDK5::::5.6:C;CDK7::::5.6:C;KPCD::::5.6:C;AURKB::::5.6:C;M4K4::::5.6:C;KPCE::::5.52:C;AKT1::::5.5:C;MYLK::::5.44:C;KPCG::::5.4:C;KS6A5::::5.3:C;SGK2::::5.2:C;AKT3::::5.2:C;CCL2::::5.16:C;CHK2::::5.1:C;IPKA|||
Sulthiame|exp|CAH2::::8.05:DC;CAN::CANAL::8.05:C;CAH9::::7.37:C;CAH15::MOUSE::7.19:C;CAH6::::6.87:C;CAH1::::6.43:C;MTCA2::MYCTU::6.18:C;CAN::YEAST::5.99:C;MTCA1::MYCTU::5.29:C|||
Parecoxib|ok|PGH2:::inh::D;TRFL|CP3A4:::sub::D;CP2C9:::inh::D||
Efaproxiral|inv|HBA;HBB|||
Triclosan|ok_inv|LMNA::::7.5:C;CBR1::::7.22:C;FABI::STAAR::7.15:DC;TAU::::6.7:C;INHA::MYCTU::6.7:DC;FABI::ECOLI::6.37:DC;FABI::BACSU::6.3:C;HS90A::::5.11:C;PGDH::::5.1:C;PERT:::inh::D;PPARG;NR1I3:::ANT::D;ANDR;NR1I2;Enoyl_acyl_carrier_protein_reductase_NADH::BACAN:::D;FABI::HELPY:::D|||
Thiamphenicol|exp_inv|STRP::STRP1::6.13:C;DRAA::ECOLX:::D|||
Dapivirine|inv|POL::HV1B1:::D|||
Diloxanide|exp||||
Ethyl_biscoumacetate|out||CP3A4:::sub::D;GLNA:::inh::D||
Azidocillin|exp|PBP2A::STRR6:inh::D;PBP1B::STRR6:inh::D;PBP3::STREE:inh::D;PBPA::STRR6:inh::D;PBP2::STRR6:inh::D||S22A5:::inh::D;S15A1:::inh::D;S15A2:::inh::D|
Pipazethate|exp||||
Salicylamide|ok|RORG::MOUSE::5.6:C;TAU::::5.05:C|||
Sulfamoxole|exp|Dihydropteroate_synthetase::PLAFA:inh::D|CP2C9:::inh::D||
Antazoline|ok|LMNA::::8.6:C;IMPA1::RAT::6.3:C;CP2D6::::5.6:C;HRH1:::ant::D|||
Chloropyramine|exp|CP2D6::::7.7:C;CP2CJ::::5.2:C;HRH1:::ant::D|||
Dimetindene|ok_inv|HRH1:::ant:9.16:DC;ACM2:::ant:7.35:DC;ACM3::::6.72:C;ACM1::::6.58:C;ACM4::::6.39:C;ACM5::::6.1:C|||
Isothipendyl|exp|HRH1:::ant::D|||
Tymazoline|exp||||
Nandrolone_decanoate|ok_ill|TAU::::5.3:C;ANDR:::ago::D|AOFA:::inh::D;AOFB:::inh::D;CP19A:::ind::D||
Roxatidine_acetate|exp|HRH2::CAVPO::7.41:C;HRH2:::ant:6.6:DC|||
Bopindolol|exp|ADRB2:::pag:7.85:DC;ADRB1:::pag:7.57:DC;5HT1A::RAT::6.82:C;ADRB3::::6.46:DC;5HT2A::::6.34:C;5HT2B::::6.01:C;5HT1B;5HT1A|CP2D6:::sub:5.26:DC||
Bupranolol|exp|ADRB3:::ant::D;ADRB2:::ant::D;ADRB1:::ant::D|CP2D6:::sub::D||
Dichloroacetic_acid|ok_inv|LMNA::::7.15:C;LEF::BACAN::5.3:C;MAAI;PDK1:::inh::D|||
Cinitapride|inv|5HT1A:::ago::D;5HT2A:::ant::D;5HT4R:::ago::D|||
Tofisopam|exp|PDE2A:::inh::D;PDE3A:::inh::D;PDE10:::inh::D;PDE4A:::inh::D|CP3A4:::inh::D||
Nadroparin|ok_inv|ANT3:::pot::D;LYAM3:::inh::D;FOS:::inh::D;MYC:::inh::D|||
Triflusal|ok_inv|CP2CJ::::5.4:C;PDE10:::ant::D;NOS2:::ago::D;NFKB1:::ant::D;PGH1:::ant::D|||ALBU:::sub::D
Lurasidone|ok_inv|DRD2:::ant::D;5HT2A:::ant::D;5HT7R:::ant::D;5HT1A:::ant::D;ADA2C:::ant::D;ADA2A|CP3A4:::sub::D||
Ticagrelor|ok|P2Y12:::inh:8.7:DC;P2Y12::RAT::5.38:C|CP2C9:::inh::D;CP2D6:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Hyaluronic_acid|ok_vet|CD44;ICAM1;HMMR;NCAN:::bin::D;CSPG2:::bin::D;C1QBP:::bin::D;HPLN1:::bin::D;HPLN3:::bin::D;HPLN4:::bin::D;HABP2:::bin::D;LAYN:::bin::D;STAB2:::bin::D;TSG6:::bin::D;IMPG2:::bin::D;HABP4:::bin::D|||
Tafluprost|ok|PF2R:::ago::D|PGH2:::ind::D||
Ivacaftor|ok|CFTR:::pot:8.52:DC;CFTR:F508del::pot:8.52:DC;CFTR:G551D::pot:6.63:DC|CP3A5:::sub::D;CP3A4:::inh::D|MDR1:::inh::D|A1AG1:::car::D;ALBU:::car::D
Azilsartan_medoxomil|ok_inv|AGTR1:::ant::D|||
Spinosad|ok_inv_vet||||
Ioflupane_I_123|ok|||SC6A3|
Deferiprone|ok|FFP::BACIU::5.85:C;KDM4E::::5.1:C|UD16:::sub::D||
Lomitapide|ok_inv|MTP:::ant:9.1:DC|CP3A4:::sub::D|MDR1:::inh::D|
Vismodegib|ok_inv|SMO::MOUSE::8.82:C;SHH::MOUSE::8.52:C;SMO:::ant:8.29:DC;SHH::::7.82:C;ALBU::RAT::5.24:C|CP2CJ:::inh::D;CP2C8:::inh::D;CP3A4:::sub::D;CP2C9:::inh::D|ABCG2:::inh::D;MDR1:::sub::D|ALBU:::sub:5.26:DC;A1AG1:::sub::D
Spaglumic_Acid|exp|FOLH1:::lig::D||S36A1:::sub::D|
Temocapril|exp_inv|ACE:::inh::D||S15A1;SO1A2|
N_methylnicotinamide|exp||AOXA:::sub::D|S22A2;S47A1:::sub::D;S47A2:::sub::D|
Acetylcarnitine|ok_inv|||S22AL::MOUSE:sub::D;S22A5|
Pitavastatin|ok|HMDH::RAT::8.39:C;ITAL;HMDH:::inh::D|CP2C8:::sub::D;CP2C9:::sub::D;UD13:::sub::D;UD2B7:::sub::D|ABCBB:::sub::D;MRP2:::sub::D;MDR1:::sub::D;ABCG2:::sub::D;NTCP:::sub::D;SO2B1:::sub::D;SO1B3:::sub::D;SO1B1:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Cholecystokinin|ok_inv|CCKAR:::ago::D;RAF1:::ago::D;MK03;EGF;KPCB:::ago::D;GASR:::ago::D||SO1B3:::sub::D;SO1B1:::inh::D;SO2B1:::inh::D|
Rilpivirine|ok|NR1I2:::ago::D;Reverse_transcriptase_RNaseH::9HIV1:inh::D|CP2D6:::inh::D;CP2B6:::inh::D;CP2CJ:::sub::D;CP3A4:::inh::D|SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|ALBU
Crizotinib|ok|MET:::inh:9.7:DC;MET:M1250T::inh:9.26:DC;ALK:::inh:9.19:DC;ROS1::::9.15:C;MET:Y1235D::inh:8.82:DC;NTRK2::::8.7:C;MERTK::::8.44:C;TIE2::::8.3:C;EPHB6::::8.22:C;UFO::::8.11:C;ALK:L1196M::inh:8.09:DC;ABL1:T315I:::8.:C;LTK::::7.92:C;SLK::::7.74:C;ABL1::::7.62:C;RON::::7.6:C;LCK::::7.52:C;IRAK3::::7.51:C;ABL1:H396P:::7.48:C;M4K1::::7.41:C;STK10::::7.36:C;IRAK1::::7.31:C;PLK4::::7.22:C;EPHA6::::7.19:C;M3K2::::7.14:C;ABL1:Y253F:::7.13:C;AURKB::::7.12:C;M4K3::::7.12:C;RON::MOUSE::7.1:C;M4K2::::7.1:C;M4K5::::7.1:C;NTRK3::::7.09:C;AURKA::::7.05:C;NTRK1::::7.02:C;ABL1:M351T:::7.01:C;ABL1:Q252H:::7.01:C;EPHA2::::7.:C;INSR::::6.99:C;TNI3K::::6.96:C;BLK::::6.96:C;M3K3::::6.96:C;TIE1::::6.96:C;NUAK2::::6.92:C;EPHB1::::6.92:C;CSKP::::6.85:C;EPHA1::::6.85:C;IGF1R::::6.84:C;ALK:F1174L::inh:6.78:DC;ABL1:E255K:::6.77:C;M3K12::::6.77:C;FAK2::::6.72:C;SIK2::::6.7:C;JAK3::::6.7:C;TYK2::::6.68:C;FLT3:D835Y:::6.68:C;CSF1R::::6.68:C;BMR1B::::6.64:C;M3K13::::6.64:C;MUSK::::6.64:C;SBK3::::6.62:C;FER::::6.57:C;EPHA8::::6.55:C;JAK2::::6.54:C;FAK1::::6.51:C;TNK1::::6.49:C;CDK7::::6.48:C;JAK1::::6.48:C;DCLK1::::6.48:C;EPHA4::::6.44:C;DCLK2::::6.43:C;TESK1::::6.42:C;CD11A::::6.38:C;ACVR1::::6.36:C;DUSTY::::6.35:C;FES::::6.35:C;TIE2::MOUSE::6.35:C;ABL2::::6.34:C;EPHA7::::6.33:C;ALK:C1156Y::inh:6.32:DC;TAOK3::::6.31:C;FLT3:D835H:::6.3:C;DDR1::::6.29:C;MK07::::6.29:C;KPCD3::::6.29:C;SRC::::6.25:C;EPHB4::::6.24:C;STK4::::6.24:C;ABL1:F317L:::6.23:C;ALK:G1269A::inh:6.22:DC;INSRR::::6.22:C;STK35::::6.21:C;ALK:S1206Y::inh:6.2:DC;KS6B1::::6.19:C;FGR::::6.17:C;LIMK2::::6.16:C;TBK1::::6.16:C;EPHA3::::6.15:C;IKKE::::6.15:C;FLT3::::6.14:C;BMP2K::::6.13:C;CD11B::::6.12:C;ACK1::::6.12:C;ANKK1::::6.11:C;YES::::6.11:C;NEK9::::6.1:C;KIT:V559D-T670I:::6.1:C;TYRO3::::6.1:C;LIMK1::::6.08:C;TXK::::6.07:C;FLT3:N841I:::6.07:C;ACV1B::::6.07:C;TAOK2::::6.05:C;RIPK2::::6.05:C;FLT3:K663Q:::6.05:C;LYN::::6.03:C;M3K19::::6.01:C;EPHA5::::6.:C;KPCD1::::6.:C;ULK1::::6.:C;TGFR1::::6.:C;STK3::::6.:C;ALK:L1152R::inh:5.99:DC;COQ8B::::5.96:C;E2AK2::::5.96:C;M3K1::::5.96:C;ABL1::MOUSE::5.94:C;ALK:G1202R::inh:5.94:DC;TAOK1::::5.92:C;RET:M918T:::5.89:C;FYN::::5.89:C;SBK1::::5.89:C;DMPK::::5.85:C;KKCC2::::5.82:C;RIPK1::::5.8:C;ULK2::::5.8:C;M3K7::::5.74:C;SRPK1::::5.74:C;ITK::::5.7:C;RET:V804L:::5.68:C;RIPK4::::5.68:C;CDKL2::::5.68:C;VGFR1::::5.64:C;AAK1::::5.64:C;AAPK1::::5.62:C;KSYK::::5.6:C;FGFR3::::5.57:C;ABL1:F317I:::5.57:C;EGFR:G719C:::5.57:C;EGFR:L861Q:::5.57:C;STK26::::5.55:C;M3K15::::5.55:C;FRK::::5.54:C;FLT3:R834Q:::5.52:C;PI51A::::5.49:C;MP2K3::::5.48:C;ROCK2::::5.48:C;FGFR3:G697C:::5.46:C;IRAK4::::5.44:C;HIPK4::::5.44:C;BMX::::5.44:C;KIT:D816V:::5.43:C;ROCK1::::5.43:C;DYRK2::::5.4:C;RIOK3::::5.4:C;GRK4::::5.38:C;ZAP70::::5.38:C;AURKC::::5.37:C;MINK1::::5.36:C;NIM1::::5.34:C;IKKB::::5.26:C;NEK7::::5.24:C;RIOK1::::5.21:C;ULK3::::5.17:C;BTK::::5.11:C;SRPK3::::5.09:C|CP3A4,CP343,CP3A5,CP3A7:::inh::D;CP2B6:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Ulipristal|ok|PRGR:::mod::D;GCR:::ant::D;ANDR|CP3A4:::sub::D;CP1A2:::sub::D||ALBU:::sub::D;A1AG1:::sub::D
Fingolimod|ok_inv|S1PR5:::mod:9.52:DC;S1PR4::::9.52:C;S1PR1::::9.52:C;S1PR3::::8.52:C;HDAC1:::inh::D|CP4FC:::sub::D;CP2E1:::sub::D;SPHK1:::sub::D;CP4F2:::sub::D||
Tesamorelin|ok_inv|GHRHR:::bin::D|||
Brentuximab_vedotin|ok_inv|TNR8:::bin::D|CP3A4:::inh::D|ABCB5:::sub::D|
Eribulin|ok_inv|TBB1;BCL2|||
Gabapentin_enacarbil|ok_inv|CA2D1;CA2D2||SC5A8:::sub::D;SC5A6:::sub::D|
Boceprevir|ok_out|CMA1::::7.49:C;CATK::::7.4:C;CATL2::::7.12:C;CATS::::6.92:C;CATL1::::6.12:C;CATF::::5.96:C;CATB::::5.21:C;Genome_polyprotein::9HEPC:inh::D|CP3A5:::inh::D;CP3A4:::inh::D|MDR1:::inh::D|
Fidaxomicin|ok|RNA_polymerase_sigma_factor_SigA::PEPD6:inh::D|CP3A4:::inh::D|MDR1:::inh::D|
Cabozantinib|ok_inv|VGFR2:::ant:10.46:DC;MET:::ant:8.89:DC;RET:::ant:8.52:DC;KIT::::8.4:C;RET:S891A::ant:8.3:DC;FLT3::::8.22:C;RET:Y791F::ant:8.15:DC;UFO::::8.15:C;FGFR1::::7.95:C;VGFR1::::7.92:C;RET:G691S::ant:7.85:DC;TIE2::::7.84:C;RET:M918T::ant:7.74:DC;RET:V804L::ant:6.64:DC;RET:V804M::ant:6.45:DC;AURKA::::5.47:C|CP2C8:::inh::D;CP2C9:::sub::D;CP3A4:::sub::D||
Taliglucerase_alfa|ok_inv|Glucocerebroside|||
Ruxolitinib|ok|JAK2:::inh:10.44:DC;JAK1:::inh:10.05:DC;TYK2::::9.4:C;JAK3::::8.7:C;M3K2::::7.39:C;KCC2A::::7.34:C;ROCK2::::7.28:C;ROCK1::::7.22:C;DCLK1::::7.17:C;DAPK1::::7.14:C;LRRK2:G2019S:::7.05:C;KCC2D::::7.05:C;DAPK3::::7.05:C;DAPK2::::7.01:C;GAK::::7.:C;KCC2G::::7.:C;KS6A1::::6.92:C;AAK1::::6.92:C;KCC1D::::6.92:C;PLK1::::6.89:C;KS6A5::::6.85:C;M3K3::::6.82:C;KS6A6::::6.82:C;KS6A2::::6.82:C;ULK2::::6.72:C;RET:V804M:::6.72:C;PLK4::::6.7:C;MKNK2::::6.7:C;BMP2K::::6.68:C;DCLK3::::6.59:C;M3K19::::6.57:C;RET:V804L:::6.55:C;LRRK2::::6.54:C;IRAK1::::6.54:C;ULK1::::6.52:C;TAOK2::::6.51:C;KCC2B::::6.51:C;NUAK2::::6.49:C;NTRK3::::6.48:C;KS6A4::::6.47:C;NTRK2::::6.44:C;MYLK::::6.44:C;ANKK1::::6.41:C;LTK::::6.36:C;CLK2::::6.34:C;MP2K3::::6.33:C;KCC1A::::6.33:C;TTK::::6.32:C;STK16::::6.31:C;KPCE::::6.28:C;MAST1::::6.28:C;GRK7::::6.27:C;TAOK3::::6.23:C;RET:M918T:::6.2:C;MARK2::::6.18:C;KGP2::::6.16:C;PLK3::::6.15:C;RK::::6.14:C;RET::::6.14:C;M3K7::::6.14:C;DCLK2::::6.12:C;DYR1A::::6.04:C;BMPR2::::6.03:C;HIPK2::::6.:C;PHKG2::::6.:C;NEK3::::5.96:C;ABL1:H396P:::5.96:C;M3K15::::5.96:C;HIPK3::::5.92:C;IKKE::::5.92:C;RIOK2::::5.92:C;HIPK1::::5.92:C;TAOK1::::5.89:C;PAK5::::5.89:C;SIK3::::5.89:C;SBK1::::5.89:C;CSKP::::5.82:C;ALK::::5.82:C;PLK2::::5.82:C;NTRK1::::5.82:C;PAK4::::5.8:C;TBK1::::5.77:C;CLK4::::5.77:C;MP2K4::::5.74:C;BMR1B::::5.74:C;KC1A::::5.74:C;MP2K1::::5.72:C;STK39::::5.72:C;RIOK3::::5.7:C;M4K2::::5.7:C;ABL1:Q252H:::5.7:C;SRPK1::::5.68:C;RIPK4::::5.68:C;BRAF::::5.66:C;ABL1:E255K:::5.66:C;ABL1:F317L:::5.66:C;MELK::::5.66:C;KCC1G::::5.66:C;IKKB::::5.64:C;ULK3::::5.62:C;RIOK1::::5.6:C;ERN1::::5.6:C;ACK1::::5.59:C;OXSR1::::5.57:C;PAK6::::5.54:C;EPHB6::::5.51:C;STK26::::5.51:C;SRPK3::::5.48:C;CDK7::::5.48:C;CSK22::::5.48:C;PI4KB::::5.47:C;ST17B::::5.46:C;DMPK::::5.46:C;DYRK2::::5.43:C;ABL1::::5.43:C;MP2K2::::5.4:C;VRK2::::5.4:C;BRAF:V600E:::5.38:C;M3K1::::5.38:C;PKNB::MYCTU::5.38:C;CSK21::::5.38:C;MK08::::5.32:C;NEK7::::5.31:C;PHKG1::::5.24:C;SBK3::::5.24:C;ST17A::::5.21:C;ABL1:M351T:::5.21:C;EPHA3::::5.21:C;GRK4::::5.21:C;STK25::::5.2:C;KIT:A829P:::5.2:C;KIT:D816H:::5.2:C;KIT:D816V:::5.15:C;AURKC::::5.06:C|CP3A4:::sub::D||
Belimumab|ok|TN13B:::neu::D|||
Teriflunomide|ok|PYRD::RAT::8.05:C;PYRD:::inh:7.52:DC;PYRD::MOUSE::7.16:C|CP1A2:::ind::D;CP2C8:::inh::D|SO1B1:::inh::D;ABCG2:::inh::D|
Vemurafenib|ok|BRAF:V600E::inh:8.4:DC;BRAF:::inh:7.7:DC;BRAF:K97R::inh:7.64:DC;RAF1::::7.32:C;VGFR2::::6.44:C;ARAF::::6.02:C;HEMH::::5.3:C|CP2B6:::ind::D;CP2C8:::inh::D;CP2C9:::inh::D;CP3A4:::sub_ind::D;CP2D6:::inh::D;CP1A2:::inh::D|ABCG2:::inh::D;MRP1:::inh::D|A1AG1:::sub::D;ALBU:::sub::D
Linagliptin|ok|DPP4:::inh:10.:DC;SEPR::::7.15:C;ACM1::::6.53:C;SEPR::MOUSE::6.43:C|CP3A4:::inh::D|S22A3:::inh::D;S22A2:::inh::D;S22A1:::inh::D;MDR1:::sub::D|
Perampanel|ok|GRIA1:::ant:6.61:DC|CP2B6:::sub_ind::D;CP1A2:::sub::D;CP3A5:::sub::D;CP3A4:::sub_ind::D||
Gadoxetic_acid|ok|||SO1B1:::sub::D;SO1B3:::sub::D;MRP3:::sub::D;MRP2:::sub::D;MRP4:::sub::D|
Aflibercept|ok|VEGFA:::bin::D;PLGF:::bin::D;VEGFB:::bin::D|||
Asparaginase_Erwinia_chrysanthemi|ok_inv||||THBG:::inh::D
Icosapent_ethyl|ok_inv_nutra||||
Ocriplasmin|ok|FINC:::cli::D;A2MG:::lig::D;A2AP:::lig::D|||
Carfilzomib|ok_inv|PSB5:::inh:8.08:DC;PSMD1::::8.07:C;PSB8:::inh:7.85:DC;PSB10:::inh::D;PSB2:::inh::D;PSB9:::inh::D;PSB1:::inh::D||MDR1:::sub::D|
Linaclotide|ok|GUC2C:::ago::D|||
Mirabegron|ok|ADRB3:::ago::D|CP3A4:::sub::D;CP2D6:::inh::D;CHLE:::sub::D|MDR1:::inh::D;SO1A2:::sub::D|ALBU:::sub::D;A1AG1:::sub::D
Peginesatide|ok_inv|EPOR:::sti::D|||
Tofacitinib|ok_inv|JAK3:::inh:9.8:DC;JAK2:::ant:9.24:DC;JAK1:::inh:9.17:DC;TYK2::::8.44:DC;DCLK3::::8.35:C;JAK3::MOUSE::7.32:C;JAK1::MOUSE::7.3:C;TNK1::::6.92:C;PKN1::::6.77:C;NUAK2::::6.62:C;ROCK2::::6.38:C;LCK::::6.34:C;ROCK1::::6.33:C;KS6A6::::6.27:C;LRRK2:G2019S:::6.26:C;KS6A2::::6.22:C;FYN::::5.96:C;PKN2::::5.92:C;KCC1A::::5.92:C;DMPK::::5.92:C;LRRK2::::5.89:C;KS6A1::::5.85:C;KCC1D::::5.8:C;MKNK2::::5.8:C;KPCD::::5.7:C;PKNB::MYCTU::5.7:C;JAK2::MOUSE::5.69:C;ABL1:T315I:::5.66:C;KCC2D::::5.57:C;RET:M918T:::5.48:C;KCC2A::::5.46:C;GRK7::::5.37:C;STK3::::5.37:C;ABL1:H396P:::5.35:C;M4K2::::5.32:C;ULK3::::5.19:C;DCLK1::::5.17:C;BMP2K::::5.15:C|CP2CJ:::sub::D;CP3A4:::sub::D||ALBU
Regorafenib|ok|HYES::::9.3:C;BRAF:::inh:7.55:DC;GLRA1::::5.74:C;RET:::inh::D;ABL1:::inh::D;FRK:::inh::D;MK11:::inh::D;RAF1:::inh::D;EPHA2:::inh::D;NTRK1:::inh::D;DDR2:::inh::D;TIE2:::inh::D;FGFR2:::inh::D;FGFR1:::inh::D;PGFRB:::inh::D;PGFRA:::inh::D;KIT:::inh::D;VGFR3:::inh::D;VGFR2:::inh::D;VGFR1:::inh::D|UD11:::inh::D;CP2B6:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;UD19:::inh::D;CP3A4:::inh::D|ABCG2:::inh::D;MDR1:::inh::D|
Aclidinium|ok|ACM3:::ant:8.36:DC;ACM5:::ant::D;ACM4:::ant::D;ACM2:::ant::D;ACM1:::ant::D|CHLE:::sub::D||
Glucarpidase|ok_inv|Methotrexate:::met::D|||
Enzalutamide|ok|ANDR:::inh:7.68:DC;ANDR::RAT::6.53:C|CP3A5:::sub_ind::D;CP2B6:::inh::D;CP2CJ:::ind::D;CP2C9:::sub_ind::D;CP3A4:::sub_ind::D;CP2C8:::inh::D|MDR1:::inh::D|THBG:::sub::D;ALBU:::sub::D
Teduglutide|ok|GLP2R::RAT::10.1:C;GLP2R:::ago:10.05:DC|||
Ponatinib|ok_inv|ABL1:::inh:10.3:DC;FLT3:::inh:9.52:DC;ABL1:T315I::inh:9.52:DC;ABL1:Q252H::inh:9.49:DC;ABL1:M351T::inh:9.39:DC;ABL1:H396P::inh:9.37:DC;ABL1:Y253F::inh:9.3:DC;FGFR1:::inh:9.15:DC;RET:::inh:9.05:DC;SRC::CHICK::9.05:C;ABL1:E255K::inh:8.97:DC;ABL1:G250E::inh:8.84:DC;VGFR2:::inh:8.77:DC;KIT:::inh:8.77:DC;SRC:::inh:8.52:DC;PGFRA:::inh::D;LYN:::inh::D;LCK:::inh::D;FGFR4:::inh::D;FGFR3:::inh::D;FGFR2:::inh::D;TIE2:::inh::D;BCR:::inh::D|CP3A5:::sub::D;CP2D6:::sub::D;CP2C8:::inh::D;CP3A4:::sub::D|ABCG2:::inh::D;MDR1:::inh::D|
Raxibacumab|ok|PAG::BACAN:abo::D|||
Bedaquiline|ok|ATPL::BACP3::6.3:C;ATPL::MYCTU:inh::D|CP3A4:::sub::D||
Certolizumab_pegol|ok|TNFA:::neu::D|AK1A1:::sub::D||
Formestane|ok_out|CP19A::::7.57:C|CP3A4:::ind::D||
Fluticasone_furoate|ok|GCR:::ago:10.4:DC;MCR:::ant::D;PRGR:::ago::D|CP2C8:::inh::D;CP3A7:::sub::D;CP3A5:::duo::D;CP3A4:::duo::D||CBG;SO1B1:::::DC;MDR1:::::DC
Canagliflozin|ok|SC5A2:::inh:8.17:DC;SC5A1::::5.72:C|CP3A4:::sub::D;UD2B4:::sub::D;UD19:::sub::D|ABCG2;MRP2:::sub::D;MDR1:::inh::D|A1AG1:::sub::D
Dimethyl_fumarate|ok_inv|KEAP1:::bin::D;TF65|||
Glycerol_phenylbutyrate|ok||LIPP:::sub::D;CP3A4:::ind::D;CP2D6:::inh::D||
Pomalidomide|ok|PGH2:::inh::D;TNFA:::inh::D;CRBN:::inh::D|CP3A4:::sub::D;CP1A2:::sub::D|MDR1:::sub::D|
Trametinib|ok|MP2K2:::ant:8.8:DC;MP2K1:::ant:8.47:DC|CP3A4:::ind::D;CP2C8:::inh::D||
Dabrafenib|ok_inv|BRAF:::ant:9.4:DC;BRAF:V600E::ant:9.:DC;ARAF::::7.59:C;RAF1:::ant:6.82:DC;TGFR1::::5.43:C;LIMK1:::ant::D;NEK11:::ant::D;SIK1:::ant::D|CP2C9:::ind::D;CP2B6:::ind::D;CP2C8:::inh::D;CP3A4:::sub_ind::D|S22A8:::inh::D;S22A6:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::sub::D|
Radium_Ra_223_Dichloride|ok_inv||||
Afatinib|ok|EGFR:G719C::inh:10.:DC;EGFR:::inh:9.96:DC;EGFR:G719S::inh:9.72:DC;EGFR:L858R::inh:9.7:DC;EGFR:L861Q::inh:9.64:DC;ERBB2:::inh:9.24:DC;EGFR:T790M::inh:9.21:DC;ERBB2:T790M::inh:9.01:DC;EGFR:L858R-T790M::inh:8.96:DC;ERBB4:::inh:8.2:DC;GAK::::7.1:C;BLK::::6.66:C;ABL1:F317L:::6.64:C;IRAK1::::6.62:C;EPHA6::::6.47:C;HIPK4::::6.44:C;ABL1:Q252H:::6.42:C;ABL1:E255K:::6.38:C;PHKG2::::6.33:C;ABL1:H396P:::6.3:C;ABL1::::6.24:C;LCK::::6.24:C;ABL1:F317I:::6.12:C;ABL1:Y253F:::6.08:C;ABL1:T315I:::6.06:C;DYR1A::::6.01:C;ABL1:M351T:::5.92:C;KC1E::::5.89:C;PHKG1::::5.89:C;MK14::::5.89:C;MP2K5::::5.89:C;FRK::::5.85:C;FLT3:D835Y:::5.85:C;MKNK2::::5.8:C;DYRK2::::5.74:C;FLT3:D835H:::5.74:C;MKNK1::::5.74:C;MK10::::5.7:C;MK09::::5.68:C;HCK::::5.66:C;MET::::5.66:C;ST17A::::5.64:C;MET:Y1235D:::5.59:C;RIPK2::::5.57:C;DYR1B::::5.55:C;SRC::::5.55:C;CTRO::::5.54:C;TXK::::5.51:C;EPHB6::::5.51:C;KS6A6::::5.51:C;SLK::::5.43:C;STK10::::5.37:C;ERBB3::::5.35:C;SBK1::::5.32:C;UFO::::5.28:C;MET:M1250T:::5.22:C;FLT3:N841I:::5.21:C||ABCG2:::inh::D;MDR1:::inh::D|
Ferric_carboxymaltose|ok||||
Levomilnacipran|ok_inv|SC6A4::RAT::8.07:C;SC6A2:::inh:7.4:DC;SC6A4:::inh:6.49:DC;SC6A3::::5.49:C;NMDZ1::RAT::5.2:C|CP2J2:::sub::D;CP2D6:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP3A4:::sub::D|MDR1:::sub::D|
Adrafinil|out||||
Arsthinol|exp||||
Dolutegravir|ok|SGMR1::CAVPO::7.15:C;Integrase::9HIV1:inh::D|UD19:::sub::D;UD13:::sub::D;CP3A4,CP343,CP3A5,CP3A7:::sub::D;UD11:::sub::D|S22A2:::inh:5.72:DC;S22A8:::inh::D;S22A6:::inh::D;ABCG2:::sub::D|MDR1:::sub::D
Riociguat|ok|GCYA2:::ago::D|CP1A1:::sub::D;CP3A4:::sub::D;CP2C8:::sub::D;CP2J2:::sub::D|ABCG2:::sub::D|ALBU:::sub::D;A1AG1:::sub::D
Macitentan|ok|EDNRA:::ant:9.3:DC;EDNRB:::ant:6.41:DC|CP2CJ:::sub::D;CP3A4:::sub::D||ALBU:::bin::D
Luliconazole|ok|CP51::CANAL:inh::D|CP2CJ:::inh::D;CP3A4:::inh::D||
Sofosbuvir|ok|POLG::HCVH::5.82:C;RNA_dependent_RNA_polymerase::9HEPC:inh::D|NDKA:::sub::D;KCY:::sub::D;HINT1:::sub::D;Q6LAP9:::sub::D;PPGB:::sub::D|ABCG2:::sub::D;MDR1:::sub::D|
Obinutuzumab|ok_inv|CD20:::abo::D|||
Chlorcyclizine|ok|HRH1:::ant::D|||
Magaldrate|ok_out||||
Letosteine|exp||||
Kebuzone|exp||||
Isoxsuprine|ok_out||||
Isoxicam|ok_out|LMNA::::6.05:C|||
Isoconazole|ok|CP17A::::6.21:C|||
Isoaminile|ok_out||||
Iotroxic_acid|exp_out||||
Iopanoic_acid|ok_out||||
Iopamidol|ok|LMNA::::5.85:C|||
Iodamide|out|LMNA::::7.5:C|||
Inositol_nicotinate|ok_out|HCAR3:::ago::D;HCAR2:::ago::D|ATPB:::inh::D;DGAT2:::inh::D|SC5A8:::sub::D|
Indoramin|out|ADA1A:::ant:8.7:DC;ADA1A::BOVIN::7.92:C;ADA1B::RAT::7.61:C;ADA1B::::7.6:C;ADA1D::::6.96:C;ADA2C::::6.32:C;ADA2B::::6.28:C;ADA1D::RAT::6.21:C;ADA2A::::5.65:C|||
Indoprofen|out|NPC1::::7.05:C;LYAG::::6.75:C;RAB9A::::6.5:C;FABPL::RAT::5.9:C;SMN::::5.9:C;NFKB2::::5.82:C;RORG::MOUSE::5.75:C;HD::::5.65:C;P53::::5.:C|||
Ifenprodil|ok_out|SGMR1::CAVPO::8.99:C;SGMR1::RAT::8.7:C;EBP::CAVPO::8.57:C;SGMR1::::8.41:C;NMDE2:::ant:8.:DC;NMDZ1:::ant:8.:DC;NMDE2::RAT::7.96:C;NMDZ1::RAT::7.14:C;ADA1B::RAT::7.:C;KCNH2::::7.:C;5HT1A::MOUSE::6.62:C;5HT2A::BOVIN::6.21:C;HRH1::::6.:C|||
Ibuproxam|out|LOX5::RAT::5.32:C;PGH2::RAT::5.:C|||
Hexoprenaline|exp_out||||
Hexetidine|ok_inv||||
Glibornuride|inv_out||CP2C9:::sub::D||
Gemeprost|ok_out|PE2R2:::ago::D;PE2R3:::ago::D|||
Fusafungine|ok_out||||
Fursultiamine|ok||||
Dimetotiazine|ok||||
Fluprednidene|exp||CP3A4:::sub_ind::D;CP3A5:::ind::D||
Fluocortolone|ok_out||CP3A5:::ind::D;CP3A4:::sub_ind::D||
Flumequine|out||CP1A2:::inh::D||
Fluclorolone_acetonide|ok_out||||
Flubendazole|exp_out|MK01::::5.:C|||
Floctafenine|ok_out||||
Fentonium|out||||
Fenspiride|exp|LMNA::::8.46:C;ACM1::RAT::5.25:C;TSHR::::5.1:C|||
Fendiline|out|CALM::BOVIN::6.3:C;CASR::::6.:C;5HT2B::::5.49:C|CP3A4:::sub::D||
Fenbufen|ok|LMNA::::6.55:C;PGH1::SHEEP::5.41:C;RAB9A::::5.25:C;PGH2::SHEEP::5.09:C;HIF1A::::5.:C|||
Etofibrate|exp||||
Etofenamate|exp|LMNA::::7.3:C;CP1A2::::6.5:C;CP2CJ::::5.:C|||THBG:::sub::D
Etilefrine|out|GALR3::::5.88:C|||
Etifoxine|inv_out||||
Etidocaine|ok|SCN1A::::5.46:C|||
Ethoheptazine|ok_out||||
Etamivan|out|BLM::::9.:C|||
Eprazinone|exp_out||||
Eperisone|inv|SGMR1::::8.77:C;ACM2::::6.08:C;ADA2B::::5.86:C;CP2D6::::5.31:C|CP3A4:::sub::D||
Ditazole|exp_out||||
Diosmin|ok_inv|AHR:::ago::D|||
Dimetacrine|exp_out|CP2D6::::5.4:C;CP1A2::::5.3:C;ACES:::ant::D|||
Dexetimide|out|ACM4::MOUSE::8.48:C|||
Cyclopentamine|out||||
Cyamemazine|exp||||
Barbexaclone|exp||||
Cloperastine|exp||||
Clobutinol|out|AL1A1::::6.82:C|||
Batroxobin|exp||||
Chlorphenoxamine|out||||
Cefaloridine|exp_out|NR1I2::::5.49:C;S22AB::::5.44:C;S15A2::RAT::5.07:C||S22A6:::sub:6.13:DC;S22A8:::inh:5.61:DC|
Articaine|ok||||
Carmofur|out|ASAH1::RAT::7.54:C;LMNA::::7.:C;CP2D6::::5.3:C;MK03::::5.21:C|||
Beclamide|exp||||
Carbazochrome|exp_out||||
Befunolol|exp|ADRB1;ADRB2|CP2D6:::sub::D||
Captodiame|exp|5HT2C:::ant::D;SGMR1:::ago::D;DRD3:::ago::D|||
Canrenoic_acid|ok_out||||
Butriptyline|ok|5HT2A:::ant::D;HRH1:::ant::D;SC6A4:::ant::D|||
Brotizolam|inv_out|PTAFR::::6.52:C|CP3A4:::sub::D||
Bromopride|inv|CP2D6::::5.3:C;AMPC::ECOLI::5.1:C;CP1A2::::5.:C;DRD2:::ant::D|||
Bromhexine|ok|SGMR1::::7.6:C;CP2D6::::6.71:C;SC6A4::::5.95:C|||
Bisacodyl|ok|LEF::BACAN::6.8:C;STAT6::::6.4:C;HIF1A::::6.3:C;GPR55::::6.04:C;OPRK::::6.01:C;TSHR::::5.9:C;LMNA::::5.85:C;SC6A3::::5.76:C;CP3A4::::5.1:C;CP2C9::::5.:C|||
Benzoctamine|exp||||
Benfluorex|inv_out|AMPC::ECOLI::6.1:C|||
Aliskiren|ok_inv|RENI:::inh:9.4:DC;RENI1::MOUSE::8.35:C;RENI::RAT::7.1:C|CP3A4:::sub::D||
Ledipasvir|ok|Nonstructural_protein_5A::9HEPC:inh::D||ABCG2:::tra::D;MDR1:::tra::D|
Cytisine|exp|ACHA4::RAT::9.91:C;ACHB2:::pag:9.64:DC;ACHA7::RAT::9.05:C;ACHA2::RAT::8.97:C;ACHA3::RAT::8.6:C;ACHA::::7.96:C;LMNA::::7.2:C;ACHA::TETCF::6.6:C;ACHB4::::6.55:C;ACHA7:::ago:5.85:DC;ACHA6:::ago::D;ACHA3:::ago::D;ACHA4:::ago::D|||
Secukinumab|ok|IL17:::ant::D|||
Vorapaxar|ok|PAR1:::ant:8.96:DC|CP2J2:::sub::D;CP3A4:::sub::D||
Miltefosine|ok_inv|LMNA::::5.45:C;AKT1::::5.02:C;MDR1|PLD1:::sub::D||
Vedolizumab|ok|ITA4:::abo::D;ITB7:::abo::D|||
Suvorexant|ok_inv|OX2R:::ant:9.46:DC;OX1R:::ant:9.26:DC;OX1R::MOUSE::8.77:C;OX2R::MOUSE::8.06:C|CP3A4:::sub::D||
Nivolumab|ok|PDCD1:::abo::D|||
Siltuximab|ok_inv|IL6:::aab::D|CP3A4:::ind::D||
Pembrolizumab|ok|PDCD1:::aab::D|||
Empagliflozin|ok|SC5A2:::ant:8.51:DC;SC5A1::::5.49:C|||
Eliglustat|ok|CEGT:::ant:7.8:DC|CP3A4:::sub::D;CP2D6:::inh::D||
Efinaconazole|ok|CP51::CANGA:inh::D|||
Tavaborole|ok_inv|SYLC::YEAST::5.73:C;Cytosolic_leucyl_tRNA_synthetase::CANAX:inh::D|||
Tedizolid_phosphate|ok||||
Albiglutide|ok|GLP1R:::ago::D|||
Dulaglutide|ok_inv|GLP1R:::ago::D|||
Metreleptin|ok|LEPR:::ago::D|||
Finafloxacin|ok_inv|GYRA::HAEIN:inh::D;PARC::HAEIN:inh::D;TOP2A:::inh::D|||
Netupitant|ok_inv|NK1R:::ant:9.02:DC|CP3A4:::inh::D;CP2D6:::sub::D;CP2C9:::sub::D;CP343:::sub::D||
Naloxegol|ok|OPRM:::ant::D|CP3A4:::sub::D;CP2D6:::inh::D;CP2CJ:::inh::D||
Ceftolozane|ok_inv|MRDA::ECOLI:inh::D;PBPC::ECOLI:inh::D;DACA,DACB,DACC,PBPA,PBPB,MRDA,FTSI::ECOLI:::D;Cell_division_protein::PSEAI:inh::D;Penicillin_binding_protein_1B::PSEAI:inh::D|||
Elosulfase_alfa|ok_inv||||
Blinatumomab|ok_inv|CD19:::act::D;CD3D:::act::D|||
Ibrutinib|ok|ERBB4::::10.:C;BTK:::inh:9.52:DC;BLK::::9.3:C;EGFR::::9.3:C;BMX::::9.1:C;LCK::::8.7:C;CSK::::8.66:C;FGR::::8.64:C;PTK6::::8.48:C;HCK::::8.43:C;YES::::8.19:C;ERBB2::::8.03:C;JAK3::::7.98:C;ITK::::7.93:C;LYN::::7.79:C;RET::::7.43:C;TEC::::7.11:C;ABL1::::7.06:C;FYN::::7.02:C;SRC::::6.58:C;FGFR2::::6.55:C;PXL2A::::6.05:C;FER::::5.09:C|CP2D6:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D||A1AG1,A1AG2:::sub::D;ALBU:::sub::D
Idelalisib|ok|PK3CD:::inh:8.7:DC;P85A::::7.6:C;PK3CG::::7.19:C;PK3CB::::6.25:C;PK3CA::::6.09:C;PRKDC::::5.17:C|CP3A7:::inh::D;CP343:::inh::D;CP3A5:::inh::D;CP3A4:::duo::D;CP2B6:::ind::D;CP2CJ:::inh::D;CP2C8:::inh::D;UD14:::inh::D;AOXA:::sub::D|SO1B3:::inh::D;SO1B1:::inh::D;MDR1:::inh::D;ABCG2:::sub::D|
Acipimox|ok_inv|HCAR2::::5.28:C|||
Amorolfine|ok_inv||||
Anthrax_immune_globulin_human|ok|PAG::BACAN:abo::D|||
Atosiban|ok_inv|V1AR:::ant:9.82:DC;OXYR::RAT::8.29:C;OXYR:::ant:7.96:DC;V1BR:::ant:7.36:DC;V2R:::ant:6.48:DC|||
Avibactam|ok|AMPC::ENTCL:inh:7.:DC;AMPC::PSEAE::6.89:C;BLE1::PSEAI:inh::D;Beta::ECOLX:inh::D;BLKPC::KLEPN:inh::D;Class::KLEPN:inh::D;BLA1::KLEPN:inh::D;BLA2::ECOLX:inh::D;BLA1::ECOLX:inh::D;Q939N4,Q9L5C7,Q840M4:::inh::D;BLAT::ECOLX:inh::D||S22A8:::sub::D;MRP2:::sub::D|
Cannabidiol|ok_inv|TRPA1::RAT::7.02:C;CAC1C::RAT::7.:C;CNR2::MOUSE::6.64:C;GPR55:::ant:6.35:DC;CNR1::RAT::5.9:C;CNR1:::ant:5.62:DC;CNR2:::ant:5.54:DC;NAAA:::inh::D;CP3A7:::inh::D;CP1A2:::inh::D;SODC:::inh::D;CATA:::inh::D;NQO1:::inh::D;CP1B1:::inh::D;I23O1:::inh::D;GPX1:::sti::D;GSHR:::sti::D;HMDH:::sti::D;CP17A:::inh::D;THIL:::inh::D;PGH2:::inh::D;PGH1:::inh::D;AA1R:::act::D;5HT3A:::ant::D;VDAC1;TRPV4:::act::D;TRPV3:::act::D;TRPV2:::act::D;TRPM8;TRPA1:::ago::D;CAC1I;CAC1H;CAC1G;TRPV1:::act::D;PPARG:::act::D;OPRM;OPRD;ACHA7;5HT2A:::ago::D;5HT1A:::ago::D;GPR18;GLRA3:::pot::D;GLRA1,GLRB:::alo::D;GLRA1;GPR12:::ANT::D|QOR;LOX15:::inh::D;LOX5:::inh::D;FAAH1:::inh::D;CP1A1:::inh::D;CP3A4:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;Arylalkylamine_N_acetyltransferase:::::DC;CP2D6:::sub::DC;CP3A5:::sub::DC|S29A1:::inh::D;ABCG2:::inh::D;MRP1:::inh::D|
Cefminox|exp||||
Ceritinib|ok|ALK:::ant:9.7:DC;ROS1::::8.7:C;INSR::::8.15:C;IGF1R::::8.1:C;TSSK1::::7.64:C;ALK:L1196M::ant:7.54:DC;FLT3::::7.22:C;FGFR2::::6.59:C;RET::::6.4:C;FGFR3::::6.37:C;LCK::::6.25:C;JAK2::::6.21:C;LYN::::6.08:C;EGFR::::6.05:C;FGFR4::::6.02:C;PGFRA::::5.94:C;ROCK2::::5.9:C;ABL1::::5.9:C;KCNH2::::5.9:C;KIT::::5.89:C;MET::::5.87:C;SRC::::5.77:C;NTRK2::::5.74:C;FGR::::5.71:C;MKNK2::::5.65:C;NTRK1::::5.56:C;KSYK::::5.52:C;ETV6::::5.49:C;BTK::::5.47:C;JAK1::::5.43:C;CDK2::::5.4:C;VGFR2::::5.38:C;CDK4::::5.33:C;JAK3::::5.1:C;ZAP70::::5.01:C|CP3A4:::inh::D;CP2C9:::inh::D|MDR1:::sub::D|
Ciprofibrate|ok_inv|PPARA::::6.05:DC;LMNA::::5.55:C;AMPC::ECOLI::5.3:C|||
Cobicistat|ok||CP3A4:::inh:6.82:DC;CP2D6:::inh:5.04:DC;CP343:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D|SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|
Corifollitropin_alfa|ok_inv|FSHR:::ago::D|||
Corticorelin_ovine_triflutate|ok|CRFR1:::lig::D|||
Vortioxetine|ok_inv|SC6A4:::inh::D;5HT3A:::ant::D;5HT7R:::ant::D;5HT1B:::pag::D;5HT1A:::ago::D;ADRB1:::lig::D;SC6A2:::inh::D|CP2D6:::sub::D;CP3A4:::sub::D;CP3A5:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP2A6:::sub::D;CP2C8:::sub::D;CP2B6:::sub::D||
Trimetazidine|ok_inv|CPT1B::RAT::5.89:C;CP1A2::::5.:C;THIK:::inh::D|||
Tibolone|ok_inv|SC6A4::::7.32:C;ANDR::RAT::7.12:C;ESR1:::duo:6.91:DC;CP2CJ::::5.52:C|ST1A1:::sub::D;3BHS2:::sub::D;3BHS1:::sub::D;STS:::inh::D||
Tasimelteon|ok_inv|MTR1A:::ago::D;MTR1B:::ago::D|CP3A4:::sub::D;CP1A2:::sub::D||
Sodium_oxybate|ok||HOT:::sub::D;SSDH:::sub::D||
Palbociclib|ok_inv|CDK4:::inh:8.7:DC;CCND1::::8.42:C;CDK6:::inh:8.05:DC;CDK2::::8.:C;CLK4::::7.7:C;JAK3::::7.2:C;DYR1B::::7.:C;ROCK2::::6.9:C;DAPK3::::6.9:C;CDK5::::6.5:C;CLK2::::6.5:C;KPCD3::::6.4:C;CDK9::::6.4:C;TAOK1::::6.3:C;DYR1A::::6.1:C;KS6A3::::6.1:C;AAPK1::::6.:C;M4K4::::5.9:C;M4K5::::5.8:C;ALK::::5.8:C;MK08::::5.8:C;CHK1::::5.6:C;MET::::5.6:C;PRKX::::5.6:C;RET::::5.6:C;LRRK2::::5.6:C;M4K2::::5.6:C;NEK2::::5.5:C;RON::::5.5:C;FLT3::::5.46:C;MK09::::5.4:C;PAK4::::5.4:C;CCNE1::::5.04:C|ST2A1:::sub::D;CP3A4:::inh::D|S22A1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|ALBU:::bin::D
Olaparib|ok|PARP1:::inh:9.62:DC;PARP2:::inh:9.55:DC;TNKS2::::8.28:C;TNKS1::::7.98:C;PARP3:::inh:7.34:DC;PARP6::::5.74:C|CP3A5:::sub::D;CP2B6:::ind::D;CP3A4:::inh::D|ABCG2:::inh::D;MDR1:::sub::D|
Edoxaban|ok|FA10:::inh:9.25:DC||MDR1:::sub::D|
Umeclidinium|ok|ACM1:::ant::D;ACM2:::ant::D;ACM3:::ant::D;ACM4:::ant::D;ACM5:::ant::D|CP2D6:::sub::D|MDR1:::sub::D|
Dinutuximab|ok_inv|Ganglioside_GD2:::inh::D|||
Lenvatinib|ok_inv|RET:::inh:8.82:DC;VGFR2:::inh:8.68:DC;VGFR3:::inh:8.28:DC;KIT:::inh::D;PGFRA:::inh::D;FGFR4:::inh::D;FGFR3:::inh::D;FGFR2:::inh::D;FGFR1:::inh::D;VGFR1:::inh::D|CP2D6:::inh::D;CP2CJ:::inh::D;CP2B6:::inh::D;CP1A2:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;AOXA:::sub::D;CP3A4:::duo::D|ABCBB:::inh::D;SO1B1:::inh::D;S22A2:::inh::D;S22A8:::inh::D;S22A6:::inh::D;ABCG2:::sub::D;MDR1:::sub::D|
Nintedanib|ok|FLT3:D835Y::inh:9.38:DC;FLT3:D835H::inh:9.15:DC;FLT3:::inh:9.15:DC;MP2K5::::8.74:C;PGFRB:::inh:8.7:DC;BMP2K::::8.66:C;FLT3:N841I::inh:8.59:DC;KIT:L576P:::8.57:C;KIT:V559D-T670I:::8.54:C;VGFR2:::inh:8.54:DC;PKNB::MYCTU::8.44:C;PGFRA:::inh:8.4:DC;M3K7::::8.39:C;FLT3:K663Q::inh:8.35:DC;NTRK1::::8.35:C;JAK1::::8.32:C;MELK::::8.31:C;VGFR3:::inh:8.3:DC;M3K19::::8.28:C;KIT::::8.24:C;LCK:::inh:8.21:DC;KIT:V559D:::8.2:C;JAK3::::8.09:C;PRP4B::::8.08:C;MERTK::::8.07:C;CLK1::::8.06:C;STK4::::8.05:C;M3K2::::8.03:C;RET:V804M:::8.02:C;RET:V804L:::8.01:C;ABL1:T315I:::8.:C;MP2K1::::8.:C;SRPK3::::7.92:C;UFO::::7.92:C;DDR1::::7.92:C;VGFR2::MOUSE::7.89:C;JAK2::::7.85:C;KGP1::::7.85:C;PI42B::::7.77:C;FLT3:R834Q::inh:7.77:DC;GRK4::::7.77:C;CLK4::::7.74:C;STK16::::7.74:C;STK11::::7.74:C;NTRK2::::7.72:C;CDK16::::7.68:C;INSRR::::7.68:C;NUAK2::::7.68:C;TTK::::7.66:C;RIOK1::::7.64:C;INSR::::7.62:C;ABL1:Q252H:::7.55:C;KIT:V559D-V654A:::7.54:C;RET:M918T:::7.52:C;ALK::::7.51:C;RET::::7.51:C;NTRK3::::7.49:C;VGFR1:::inh:7.47:DC;M3K3::::7.47:C;M4K1::::7.46:C;RIOK3::::7.44:C;SRPK2::::7.44:C;SRPK1::::7.43:C;TYK2::::7.43:C;ABL1:Y253F:::7.43:C;FGFR2:::inh:7.43:DC;LRRK2:G2019S:::7.43:C;FGFR1:::inh:7.42:DC;STK3::::7.42:C;MP2K2::::7.38:C;DDR2::::7.38:C;ABL1:H396P:::7.35:C;LRRK2::::7.34:C;KIT:D816V:::7.33:C;CSF1R::::7.32:C;STK26::::7.31:C;PI51A::::7.31:C;SLK::::7.29:C;ABL1:M351T:::7.28:C;PLK4::::7.28:C;TNIK::::7.28:C;BMPR2::::7.25:C;KS6A2::::7.24:C;ULK3::::7.22:C;IGF1R::::7.21:C;ABL1:E255K:::7.2:C;AAK1::::7.2:C;KS6A3::::7.19:C;ABL1::::7.19:C;FER::::7.14:C;YES::::7.1:C;FAK2::::7.09:C;MINK1::::7.09:C;AAPK2::::7.08:C;GSK3B::::7.08:C;STK10::::7.06:C;AAPK1::::7.06:C;KIT:A829P:::7.06:C;CDK17::::7.03:C;FGFR3:::inh:7.03:DC;STK24::::6.96:C;ST17A::::6.96:C;MYLK3::::6.96:C;SBK1::::6.96:C;IRAK1::::6.92:C;EPHB6::::6.85:C;M3K13::::6.85:C;PHKG1::::6.85:C;M3K12::::6.85:C;FGFR3:G697C::inh:6.85:DC;TBK1::::6.82:C;LTK::::6.82:C;M4K4::::6.82:C;SRC:::inh:6.81:DC;NUAK1::::6.8:C;CDK4::::6.8:C;IKKE::::6.77:C;KS6A1::::6.74:C;KS6B1::::6.72:C;AURKC::::6.72:C;LYN:::inh:6.71:DC;KS6A5::::6.7:C;MET::::6.7:C;TNK1::::6.68:C;ITK::::6.68:C;FAK1::::6.68:C;PAK3::::6.68:C;M3K9::::6.66:C;KS6A6::::6.64:C;KC1E::::6.64:C;RIPK1::::6.62:C;KCC1G::::6.59:C;PHKG2::::6.59:C;MK10::::6.57:C;SIK2::::6.55:C;M4K3::::6.54:C;M4K2::::6.54:C;MYLK::::6.54:C;CHK1::::6.54:C;FGR::::6.52:C;CDK7::::6.52:C;BTK::::6.51:C;KIT:D816H:::6.51:C;ULK1::::6.47:C;MET:M1250T:::6.47:C;LATS2::::6.42:C;ULK2::::6.42:C;BLK::::6.42:C;M4K5::::6.41:C;LATS1::::6.38:C;AURKB::::6.38:C;GSK3A::::6.37:C;RIPK4::::6.36:C;MYLK4::::6.36:C;MET:Y1235D:::6.34:C;CDK14::::6.33:C;CDK18::::6.29:C;STK39::::6.28:C;DCLK1::::6.27:C;EPHB1::::6.26:C;MUSK::::6.23:C;ACVR1::::6.22:C;FGFR4::::6.21:C;KS6A4::::6.21:C;KKCC1::::6.2:C;FYN::::6.2:C;MK08::::6.2:C;ABL1:F317L:::6.19:C;KPCD3::::6.19:C;ST17B::::6.17:C;SIK1::::6.17:C;M3K11::::6.15:C;KPCD2::::6.14:C;PKN1::::6.13:C;CLK2::::6.12:C;DCLK3::::6.11:C;MARK3::::6.11:C;HIPK2::::6.1:C;IRAK4::::6.09:C;STK35::::6.09:C;TXK::::6.07:C;HIPK3::::6.07:C;CSK22::::6.05:C;KKCC2::::6.04:C;EPHA6::::6.03:C;SGK3::::6.:C;KPCD1::::6.:C;RK::::6.:C;EPHB4::::5.96:C;STK33::::5.96:C;EPHA1::::5.92:C;CDPK1::PLAF7::5.92:C;FES::::5.92:C;GRK7::::5.92:C;HIPK4::::5.92:C;CDKL2::::5.89:C;OXSR1::::5.89:C;PAK5::::5.89:C;HIPK1::::5.89:C;KC1D::::5.89:C;PKN2::::5.85:C;MARK2::::5.85:C;MARK1::::5.85:C;TIE2::::5.85:C;M3K15::::5.85:C;CDK2::::5.85:C;DYR1B::::5.8:C;ACK1::::5.8:C;ICK::::5.77:C;ABL2::::5.7:C;MARK4::::5.7:C;SBK3::::5.7:C;E2AK4::::5.7:C;ERN1::::5.7:C;DAPK3::::5.68:C;MP2K3::::5.68:C;TIE1::::5.66:C;KCC1D::::5.66:C;M3K10::::5.64:C;MK07::::5.6:C;ABL1:F317I:::5.59:C;MYO3B::::5.57:C;FRK::::5.57:C;PDPK1::::5.55:C;WEE1::::5.54:C;EPHA2::::5.54:C;PAK4::::5.52:C;DAPK2::::5.49:C;PAK2::::5.48:C;ZAP70::::5.46:C;KCC2A::::5.44:C;MP2K4::::5.43:C;KCC4::::5.43:C;ROS1::::5.43:C;MYLK2::::5.4:C;TGFR1::::5.38:C;ACVL1::::5.38:C;IKKA::::5.35:C;MAST1::::5.34:C;ACV1B::::5.31:C;TYRO3::::5.31:C;IRAK3::::5.28:C;HCK::::5.28:C;KPCT::::5.26:C;KCC1A::::5.23:C;TSSK1::::5.21:C;CSK21::::5.12:C;EPHA3::::5.07:C|CP3A4:::sub::D;UD110:::sub::D;UD18:::sub::D;UD17:::sub::D;UD11:::sub::D|ABCG2;S22A1:::inh::D;MDR1:::inh::D|ALBU:::sub::D
Olodaterol|ok|ADRB2:::ago::D|CP2C9:::sub::D;CP2C8:::sub::D||
Idebenone|ok_inv|CP2CJ::::6.1:C;CP2D6::::5.52:C;CP2C9::::5.3:C;CP3A4::::5.15:C|||
Vilanterol|ok|ADRB2:::ago::D|CP3A4:::sub::D||
Ivabradine|ok|HCN4::::5.37:C;HCN1::MOUSE::5.35:C;HCN2::MOUSE::5.34:C;HCN2:::inh::D|CP3A4:::sub::D||
Benzydamine|ok|GCYB1::::5.99:C;CP1A2::::5.3:C;CP2D6::::5.1:C|||
Tetracaine|ok_vet|SCN9A::::7.25:C;AOFA::::6.5:C;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A:::inh:6.4,,,6.31,6.13,,6.28,,6.28,7.25:DC;SCN1A::::6.4:C;SCN2A::::6.31:C;SCN8A::::6.28:C;SCN5A::::6.28:C;SGMR1::::6.15:C;SCN3A::::6.13:C;5HT2A::::6.01:C;5HT2C::::5.77:C;SCN2A::RAT::5.22:C;CNGA1::BOVIN::5.17:C;RYR2:::mod::D;RYR1:::mod::D|||
Eugenol|ok|CP3A4::::5.4:C;TRPV3;ANDR:::ant::D;ESR2;ESR1|||
Potassium_alum|ok||||ALBU:::bin::D
Amylocaine|ok_out|SCN1A:::inh::D|||
Trimebutine|ok|OPRM:::ago::D;CAC1C:::inh::D;KCMA1:::inh::D;CAC1G:::act::D;ACM1:::ant::D;ACM2:::ant::D;ACM3:::ant::D;ACM4:::ant::D|CP3A4:::sub::D||
Pinaverium|ok|CAC1C::::5.76:C;CAC1S:::ant::D|CP3A4:::sub::D||
Tixocortol|ok_out|GCR:::bin::D;HDAC2:::sti::D|||
Xanthinol|ok_out|RL3:::bin::D;NNTM:::cof::D;G3P:::cof::D;IDH3A:::cof::D;ODO1:::cof::D;MDHM:::cof::D|||
Chlortetracycline|ok_inv_vet|RS7::ECOLI:inh::D;RS14::ECOLI:inh::D;RS19::ECOLI:inh::D;RS8::ECOLI:inh::D;RS3::ECOLI:inh::D;16S_ribosomal_RNA::Gut_flora:inh::D|||ALBU
Podophyllin|ok||||
Difluocortolone|ok_out|GCR:::bin::D;ANXA3:::ind::D|CP3A5:::ind::D;CP3A4:::sub_ind::D||
Benzoyl_peroxide|ok|LMNA::::8.2:C|||
Quinagolide|ok_inv|DRD1::BOVIN::7.72:C;5HT3A::RAT::5.64:C;ADA2C::RAT::5.25:C;ADA1B::RAT::5.22:C;DRD1,DRD5:::ago::D;DRD2:::ago::D|||
Somatrem|ok_out|GHR:::ago::D;IGF1R|||
Somatostatin|ok_inv|SSR1:::ago::D;SSR2:::ago::D;SSR3:::ago::D;SSR4:::ago::D;SSR5:::ago::D|CP3A4:::inh::D|MDR1:::sub::D|
Thyroid_porcine|ok||||
Elvitegravir|ok|Integrase::9HIV1:inh::D|UD14:::sub::D;CP3A4:::inh::D||
Daclatasvir|ok_inv|Nonstructural_protein_5A::9HEPC:inh::D|CP3A4:::sub:5.14:DC;CP3A7:::sub::D;CP343:::sub::D;CP3A5:::sub::D|ABCG2:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;MDR1:::inh::D|
Ancestim|ok_out|KIT:::ago::D|||
Magnesium_hydroxide|ok_inv||||
Asfotase_alfa|ok_inv|S1PR1:::ago::D;Pyrophosphate::UNK:lig::D|||
Hydroxyethyl_Starch|ok||||
Methoxy_polyethylene_glycol_epoetin_beta|ok|EPOR:::sti::D|||
Simoctocog_alfa|ok|VWF:::bin::D|||
Turoctocog_alfa|ok_inv|FA9:::act::D;FA10:::act::D;THRB:::bin::D|||
Coenzyme_M|ok_inv||GSHR:::sub::D||
Pentastarch|ok_inv||||
Nitrous_acid|ok_inv|MYG:::oxi::D;HBB:::oxi::D;HBA:::oxi::D|||
Poractant_alfa|ok||||
Colfosceril_palmitate|ok_out|AMPC::ECOLI::6.45:C|||
Diiodohydroxyquinoline|ok|HIF1A::::6.7:C;MK01::::6.53:C;RORG::MOUSE::6.45:C;MK14::::6.44:C;HS90A::::6.41:C;AA3R::::6.28:C;ACE::RABIT::6.04:C;FYN::::5.8:C;EGFR::::5.72:C;LCK::::5.61:C;AMPC::ECOLI::5.4:C;PAX8::::5.31:C;MK03::::5.28:C;COMT::RAT::5.25:C;CYSP::TRYCR::5.2:C;P53::::5.1:C;ERBB2::::5.07:C|||
Calcium_carbimide|ok_out|AL3B2:::ant::D|CATA:::sub::D||
Paraldehyde|ok_inv|LMNA::::5.:C|ALDH2:::sub::D||
Stiripentol|ok|LDHB:::inh::D;LDHA:::inh::D;GABAR:::ago::D|CP2C9:::inh::D;CP1A2:::inh::D;CP3A4:::inh::D;CP2D6:::inh::D;CP2CJ:::inh::D||
Eslicarbazepine_acetate|ok|P2RX4:::ant::D|UD11:::sub::D;CP3A4:::ind::D;CP2CJ:::inh::D||
Zucapsaicin|ok_inv|AL1A1::::5.45:C;CP3A4::::5.4:C;CP2D6::::5.2:C;LEF::BACAN::5.2:C;TRPV1:::ago::D|CP2C9:::inh:6.5:DC;CP1A2:::inh:5.8:DC;CP2CJ:::inh:5.2:DC;CP2E1:::inh::D||
Aurothioglucose|ok_out|ADCY1;ADCY2;ADCY5|||
Peginterferon_beta_1a|ok||CP1A2:::inh::D||
Dienogest|ok|PRGR:::ago::D;ANDR:::ant::D|CP3A4:::sub::D||
Medrogestone|ok|PRGR:::lig::D|CP3A4:::sub::D||ALBU:::bin::D;SHBG:::bin::D;CBG:::bin::D
Potassium_citrate|ok_inv_vet||||
Chorionic_Gonadotropin_Human|ok_vet|LSHR:::lig::D|||
Brexpiprazole|ok_inv|DRD2::RAT::9.7:C;5HT2A::RAT::8.64:C;ADA1B:::ant::D;ADA2C:::ant::D;5HT2A:::ant::D;DRD2:::ago::D;5HT1A:::ago::D|CP3A4:::sub::D;CP2D6:::sub::D||
Chromic_chloride|ok|INSR:::act::D|||
Copper|ok_inv|A4:::agi::D;SAHH:::alo::D;H2B1C;G3P;NDKA;H14;PRDX1;S10A8;RSSA;ACTG;ENOA;EF1A1;K2C8;PDIA1;PDIA3;CH60;HSP13;BIP;ENPL;TRFE;LYAR::MOUSE:::D;RS2;SRSF1;ROA2;HNRH1;HNRH3;CBID::TREDE:::D;HNRPL;SFPQ;SF3A2;RACK1;ACTN1;ACY1;ANXA4;ANXA5;CALR;KPYM;AK1A1;NB5R3;GSHR;TKT;PRDX2;PRDX6;PPIA;HSP7C;HS90A;TEBP;STIP1;Translation_elongation_factor_1_alpha_1_like_14;IF6;IF4A1;G6PI;LDHA;PGK1;TBA3D;TBB5;COF1;1433B;AATC;GSHB;HDGF;IDH3A;CLIC1;PSME1;PEBP1;PGAM1;RANG;UGDH;B2MG;SCO1;APRIO;GLRA1;HD;NEIL1;NEIL2;HPHL1:::cof::D;PAI1;S10A2;S10A4;SYUA;BDNF:::cof::D;PARK7;IAPP;TKNK;A1BG;AFAM;ANGT;FETUA;SAMP;APOA1;APOA2;APOA4;APOBR;APOC2;APOC3;APOD;APOE;APOH;ZA2G;C1QC;C1S;CO3;CO4B;C4BPA;CO5;CO8B;CO9;CFAH;CFAI;TETN;CLUS;THRB;C1QBP;GELS;HBA;HBB;CBX5;HPTR;ALS;IGHG1;IGHG4;KV320;IGLL1;ITIH2;KNG1;K2C1;K1C10;K22E;K1C9;A2GL;LUM;PGRP2;PLMN;PON1;CXCL7;A1AT;KAIN;CBG;THBG;ANT3;HEP2;PEDF;A2AP;IC1;TTHY;VTNC;APLP1:::cof::D|SODC:::cof::D;AOC1:::cof::D;LYOX:::cof::D;COX1:::cof::D;TYRO:::cof::D;DOPO:::cof::D;AMD:::cof::D;AOFA:::cof::D;ANGI:::cof::D;PRIO:::cof::D|COPT1:::sub::D;NRAM2:::sub::D;ATP7A:::sub::D;ATP7B:::sub::D;COPT2|ALBU:::bin::D;A2MG:::bin::D;CERU:::bin::D;ATOX1:::bin::D;CCS:::bin::D;COX17:::bin::D;HEPH:::bin::D;FA5:::bin::D;FA8:::bin::D;MTF1:::bin::D
Cupric_Chloride|ok_inv|PROC;CYTB|||
Gadoteric_acid|ok||||
Iothalamic_acid|ok||||
Ioversol|ok||||
Ioxilan|ok||||
Isosulfan_blue|ok||||
Technetium_Tc_99m_mebrofenin|ok|||SO1B1:::sub::D;SO1B3:::sub::D|
Technetium_Tc_99m_medronate|ok||||
Technetium_Tc_99m_oxidronate|ok||||ALBU:::bin::D
Oxygen|ok_vet|COX1:::ago::D;NOX1:::ago::D;HBA;HBB|||
Protamine_sulfate|ok|FA10;ANT3|||
Sincalide|ok|GASR::::10.3:C;CCKAR::RAT::10.05:C;CCKAR::::10.:C;CCKAR::CAVPO::9.55:C;CCKAR::MOUSE::9.52:C;GASR::MOUSE::9.52:C;GASR::RAT::9.39:C||SO1B3:::sub::D|
Sonidegib|ok_inv|SHH::MOUSE::8.26:C;SMO:::ant:8.22:DC|CP3A4:::sub::D||
Uridine_triacetate|ok_inv||||
Water|ok||||
Iron_sucrose|ok|HBA|||TRFE:::car::D
Florbetaben_18F|ok|A4:::bin:8.65:DC|CP4F2:::sub::D;CP2J2:::sub::D||
Florbetapir_18F|ok_inv|A4:::bin:8.54:DC|||
Flutemetamol_18F|ok_inv|A4:::bin::D|||
Nitrogen|ok_vet||||
Sodium_chloride|ok_vet||||
Sodium_citrate|ok_inv|CAH4::::7.:C||TXTP:::sub::D;S13A5:::sub::D;S13A2:::sub::D;ODC:::sub::D|
Helium|ok_inv_vet||||
Iopromide|ok||||
Carbon_dioxide|ok_inv_vet||||
Trypan_blue_free_acid|ok|PTN1::::5.41:C;PTP1::YEAST::5.13:C|||
Technetium_Tc_99m_tetrofosmin|ok||||MDR1:::bin::D
Technetium_Tc_99m_sestamibi|ok_inv|||MDR1:::sub::D;MRP1:::sub::D|
Technetium_Tc_99m_exametazime|ok||||
Technetium_Tc_99m_disofenin|ok||||
Technetium_Tc_99m_pyrophosphate|ok|Hydroxyapatite:::lig::D;Amorphous_calcium_phosphate:::lig::D|||
Etizolam|exp|PTAFR:::ant::D;GBRG2:::ago::D;GBRA3:::ago::D;GBRA2:::ago::D;GBRA1:::ago::D|CP2CJ:::sub::D;CP2CI:::sub::D;CP3A4:::sub::D||
Dosulepin|ok|SC6A4:::inh::D;SC6A2:::inh::D;ADA1A,ADA1B,ADA1D:::ant::D;ADA2A,ADA2B,ADA2C:::ant::D;ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D;HRH1:::ant::D;5HT2A:::ant::D;5HT1A:::ant::D|CP2D6:::inh:5.1:DC;CP2C9:::inh::D;CP2CJ:::inh::D;CP1A2:::inh::D||
Dasabuvir|ok|Nonstructural_protein_5b::9HEPC:inh::D|UD14:::inh::D;CP2D6:::sub::D;CP3A4:::sub::D;CP2C8:::sub::D|MDR1:::sub::D;ABCB5:::sub::D;ABCG2:::inh::D|
Viloxazine|ok_out|SC6A2:::inh:6.81:DC;SC6A3::::6.81:C|CP1A2:::inh::D||
Etoperidone|out|ADA1A:::ant::D;ADA2A:::ant::D;DRD2:::ant::D;ACM1:::ant::D;5HT2A:::ant::D;5HT2C:::ago::D||SC6A4:::inh::D;SC6A2:::inh::D;SC6A3:::inh::D|
Lorpiprazole|ok|5HT2A:::ant::D;5HT2C:::ant::D;ADA1A:::ant::D;ADA2A:::ant::D;HRH1:::ant::D;SC6A4:::ant::D|CP2D6:::sub::D;CP3A4:::sub::D||ALBU:::sub::D
Synephrine|exp|BLM::::8.55:C;SMN::::6.15:C;ACM1::RAT::5.85:C;NMUR2::::5.18:C;TPO::::5.:C;ADA1A,ADA1B,ADA1D|||
Moxisylyte|ok_inv|KPYM::::7.9:C;ADA1A,ADA1B,ADA1D,ADA2A,ADA2B,ADA2C:::ant:7.5,,,,,:DC;ADA1A::::7.5:C;CP1A2::::5.5:C;ACM1::RAT::5.1:C;CP2D6::::5.:C|CP3A4,CP343,CP3A5,CP3A7:::sub::D;CHLE:::sub::D||
Trimazosin|exp||||
Pegloticase|ok_inv|Uric_acid:::met::D|||
Pholcodine|ok_ill|OPRM:::ant::D;OPRK:::ant::D;OPRD:::ant::D|||
Piracetam|ok_inv|AMPC::ECOLI::5.8:C|||
Loxoprofen|ok|PGH1:::ant:5.19:DC;PGH2:::ant::D|UD2B7:::sub::D;CP3A4,CP343,CP3A5,CP3A7:::sub::D;CBR1:::sub::D||
Dexibuprofen|ok_inv|BLM::::8.55:C;PGH1:::inh:7.01:DC;CXCR2::::7.:C;END4::ECOLI::6.6:C;PGH2:::inh:6.14:DC;PGH1::SHEEP::5.83:C;PGH2::SHEEP::5.82:C;TSHR::::5.6:C;LMNA::::5.6:C;S10A7;GP1BA;PPARA;S15A1;CFTR:::inh::D;PPARG:::act::D;FABPI:::bin::D;TPA:::mod::D;TRBM:::mod::D;BCL2:::neg::D|UD2B7:::sub::D;D6RB81:::sub::D;CP2CJ:::sub::D;UD2B4:::sub::D;UD19:::sub::D;UD13:::sub::D;UD11:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D|MDR1;SO2B1;S22AB;S22A8;S22A6;SO1A2;MRP1;MRP4|ALBU
Dexketoprofen|ok_inv|CXCR2::::7.3:C|PGH1:::inh:8.72:DC;PGH2:::inh:7.57:DC||
Droxicam|out|PGH2:::inh::D;PGH1:::inh::D|||
Tolfenamic_acid|ok_inv|AK1C3::::8.1:C;TTHY::::6.82:C;CP2C9::::5.5:C;CP1A2::::5.5:C;LMNA::::5.15:C;PA21B::::5.11:C;ATG4B::::5.09:C;TAU::::5.:C;HIF1A::::5.:C;UBP2::::5.:C;PGH2:::ant::D;PGH1:::ant::D|CP3A4:::sub::D||
Bisoxatin|ok||||
Nicorandil|ok_inv|CP2C9::::5.7:C;CP2CJ::::5.4:C;ABCC9:::act::D|||
Fibrinogen_human|ok||||
Melperone|inv|DRD2:::ant::D|CP2D6:::inh::D||
Zotepine|ok_out|5HT2A:::ant:9.3:DC;HRH1::::9.21:C;5HT2C::::8.54:C;ADA1A::::8.47:C;DRD3::::8.19:C;DRD2:::ant:7.96:DC;DRD1,DRD5:::ant:7.54,:DC;DRD1::::7.54:C;DRD4::::7.41:C;ADA2A::::6.74:C;5HT1A::::6.48:C;ACM4::::6.26:C;SC6A4:::ant::D;SC6A2:::ant::D;5HT7R:::ant::D;5HT6R:::ant::D|CP3A4:::sub::D;CP1A2:::sub::D||
Barnidipine|exp|CAC1C:::ant:5.92:DC;MDR1::::5.07:C|CP3A4:::inh::D||
Conestat_alfa|ok_inv|C1R:::inh::D;C1S:::inh::D;KLKB1:::inh::D;FA12:::inh::D;THRB:::inh::D;FA11:::inh::D;TPA:::inh::D|||
Benidipine|exp|MDR1::::5.3:C;CAC1G,CAC1H,CAC1I:::ant::D;CAC1B:::ant::D;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1A:::ant::D|CP3A5:::sub::D;CP3A4:::inh::D||
Cilnidipine|inv|CAC1C::RAT::8.96:C;CAC1B:::ant:5.8:DC;MEN1::::5.75:C;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1A:::ant:5.28,,,,,,,,:DC;CAC1C::::5.28:C|CP3A4:::sub::D||
Lacidipine|ok_inv|THAS::::5.77:C;CP2CJ::::5.7:C;CP2C9::::5.7:C;DRD3::::5.68:C;AA3R::::5.64:C;ANDR::RAT::5.58:C;SC6A2::::5.25:C;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1A:::ant::D|CP3A4:::sub:6.05:DC||A1AG1:::bin::D;ALBU:::bin::D
Levamlodipine|ok_inv|CAC1C:::ant::D;CAC1D:::ant::D;NOS3:::ago::D;NOS2:::ago::D|CP3A4:::sub::D;NOS2:::ind::D;NOS3:::ind::D|MDR1:::sub::D;NTCP2:::inh::D;S22A5:::inh::D|ALBU:::bin::D
Manidipine|ok_inv|MDR1::::5.34:C;CYSP::TRYCR::5.22:C;CAC1G,CAC1H,CAC1I:::inh::D;CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1A:::inh::D|CP3A4:::inh::D;CP2CJ:::inh::D;CP2B6:::inh::D;CP1A1:::inh::D;CP2D6:::inh::D;CP2C9:::inh::D||
Methylene_blue|ok_inv|PPARG::::6.13:C;RAD52::::6.03:C;TAU::::5.9:C;NPSR1::::5.8:C;CASP6::::5.8:C;GSHR::PLAF7::5.19:C;MK01::::5.15:C;NOS1:::ant::D;GCYA2:::ant::D|||
Moxonidine|ok_inv|NISCH:::ago:8.38:DC;ADA2A:::ago:7.12:DC;NISCH::RAT::7.11:C;LMNA::::6.4:C;5HT1A::RAT::6.4:C;ADA2B::RAT::6.:C;ADA2C::::5.7:C|||
Toloxatone|exp|AOFA::BOVIN::6.42:C;AOFA::RAT::6.42:C|AOFA:::inh:5.82:DC||
Iproclozide|out||||
Dextran|ok_inv_vet||||
Tegafur|ok_inv|AMPC::ECOLI::5.8:C;RORG::MOUSE::5.3:C;TAU::::5.1:C;TYSY:::inh::D|CP3A5:::sub::D;CP2E1:::sub::D;CP2A6:::sub::D;CP2C8:::sub::D;CP1A2:::sub::D||THBG:::ind::D
Gimeracil|ok|DPYD:::inh::D|||
Bemiparin|ok_inv|FA10:::ant::D;ANT3:::ant::D;HEP2:::ant::D|||
Reviparin|ok_inv||||
Parnaparin|ok_inv||||
Certoparin|ok_inv||||
Patiromer|ok_inv|Potassium:::bin::D|||
Idarucizumab|ok||||
Lixisenatide|ok|GLP1R:::ago::D|||
Technetium_Tc_99m_tilmanocept|ok_inv|MRC1:::lig::D|||
Strontium_ranelate|ok_out||||
Picosulfuric_acid|ok||Arylsulfate_sulfotransferase_AssT::ECOK1:sub::D||
Phenylacetic_acid|ok||EST1:::sub::D||
Ubidecarenone|ok_inv_nutra|LMNA::::7.95:C;SDHA:::cof::D;NDUV3:::cof::D|HMDH:::sub::D|MDR1:::sub::D|VLDLR:::sub::D;LDLR:::sub::D
Cimetropium|exp_inv||||
Eluxadoline|ok_inv|OPRM::RAT::9.05:C;OPRM:::ago:9.:DC;OPRD::RAT::8.89:C;OPRK::CAVPO::7.26:C;OPRK:::ago::D;OPRD:::ant::D||S22A8:::sub::D;MRP2:::sub::D;SO1B1:::inh::D|
Doxofylline|exp|ADRB2:::ago::D;AA2AR:::ant::D;Phosphodiesterase_2A_cGMP_stimulated:::inh::D|CP1A2:::sub::D||
Artesunate|ok_inv|EXP1::PLAFA:inh::D|CP3A4:::sub::D;CP2A6:::sub::D||
Bismuth_subcitrate_potassium|ok_inv|CLPX::HELPY:ant::D|||
Sodium_aurothiomalate|ok_inv||UD11:::inh::D||
Choline_C_11|ok_inv||||
Activated_charcoal|ok||||
Fimasartan|inv|AGTR1::RABIT::9.38:C;AGTR1:::ant::D||ABCG2:::sub::D;SO1B1:::sub::D|
Lumacaftor|ok|CFTR:::mod:5.59:DC|CP2CJ:::ind::D;CP2C9:::duo::D;CP2C8:::duo::D;CP2B6:::ind::D;CP3A4:::ind::D|MDR1:::duo::D|ALBU:::car::D
Magnesium_trisilicate|ok||||
Molsidomine|ok_inv|THB::::7.9:C;HIF1A::::6.5:C;CP3A4::::5.9:C;LMNA::::5.2:C;ACM1::RAT::5.1:C;TYDP1::::5.05:C;END4::ECOLI::5.:C|PDE5A:::sub::D;GCYA2:::ind::DC||
Trapidil|exp|LMNA::::7.5:C;CP1A2::::5.4:C;MK01::::5.15:C;PDE1A,PDE1B,PDE1C,PDE10,PDE4A,PDE4B,PDE4C,PDE4D,PDE7B,PDE2A,PDE3A,PDE3B,PDE5A,PDE6C,PDE11,PDE7A,PDE8A,PDE8B,PDE9A,PDE6A,PDE6B:::inh::D;PGFRB:::ant::D|||
Imolamine|inv||||
Morniflumate|exp|TA2R;LT4R1:::ant::D|UD19:::inh::D;PGH2:::inh::DC;LOX5:::inh::DC||
Pipamperone|inv|ADA2A:::ant::D;5HT2B;DRD3;DRD1:::ant::D;DRD4:::ant::D;ADA1A,ADA1B,ADA1D:::ant::D;5HT2A:::ago::D;DRD2:::ant::D|||
Polyethylene_glycol|ok_vet||||
Propacetamol|exp|CNR1:::ant::D;TRPV1:::ant::D;PGH2:::ant::D;PGH1:::ant::D|CP3A4:::sub_ind::D;CP2C9:::sub::D;ARY2:::inh::D;ST2A1:::sub::D;ST1E1:::sub::D;ST1A3:::sub::D;ST1A1:::sub::D;UD110:::sub::D;UDB15:::sub::D;UD19:::sub::D;UD16:::sub::D;UD11:::sub::D;CP2D6:::sub::D;CP1A2:::sub::D;CP2E1:::sub::D;CHLE:::sub::D||
Tianeptine|inv|DRD3:::ago::D;5HT1A:::inh::D;OPRM:::ago::D;GRIA1:::mod::D|CP3A4:::sub::D||
Rolapitant|ok_inv|NK1R:::ant::D|CP2D6:::inh::D;CP3A4:::sub::D|ABCG2:::inh::D;MDR1:::inh::D|
Sacubitril|ok|NEP:::ant::D||SO1B1:::inh::D;SO1B3:::inh::D|
Iodide_I_131|ok_inv||||
Ombitasvir|ok_inv|Nonstructural_protein_5A::9HEPC:inh::D|CP2C8:::sub::D|ABCG2:::sub::D;UD14:::inh::D;MDR1:::sub::D|
Paritaprevir|ok_inv|Genome_polyprotein::9HEPC:inh::D|CP3A4:::sub::D;CP3A5:::sub::D;UD11:::inh::D|ABCG2:::inh::D;MDR1:::sub::D;SO1B1:::inh::D;SO1B3:::inh::D|
Tenofovir_alafenamide|ok|DNA_polymerase::HHV21:inh::D;Reverse_transcriptase::HBV:inh::D;Reverse_transcriptase_RNaseH::9HIV1:inh::D|NDKB:::sub::D;NDKA:::sub::D;KAD2:::sub::D;KAD1:::sub::D;CP3A4:::sub::D;EST1:::sub::D;PPGB:::sub::D|SO1B3:::sub::D;SO1B1:::sub::D;ABCG2:::sub::D;S22A8:::sub::D;S22A6:::sub::D;MRP4:::sub::D;MDR1:::sub::D|ALBU:::bin::D
Butylscopolamine|ok_inv_vet|ACM3:::ant::D;ACM2:::ant::D|||
Chondroitin_sulfate|ok_inv_nutra|BDNF;GDNF;VEGFA;CCL2|BGLR:::sub::D;HEXB:::sub::D;GALNS:::sub::D;IDS:::sub::D;IDUA:::sub::D;ARSB:::sub::D||
Alirocumab|ok|PCSK9:::inh::D|||
Evolocumab|ok||PCSK9:::inh::D||
Solithromycin|inv||CP3A4:::inh::D||
Catridecacog|ok|F13B|||
Antilymphocyte_immunoglobulin_horse|ok_inv||||
Ioxaglic_acid|ok_inv|AMPC::ECOLI::6.2:C|||
Technetium_Tc_99m_pertechnetate|ok_inv||||
Xenon_133|ok||||
Thallous_Chloride|ok||||
Synthetic_Conjugated_Estrogens_A|ok|ESR1:::lig::D|CP3A4:::sub::D||THBG:::ind::D
Synthetic_Conjugated_Estrogens_B|ok|ESR1:::lig::D|CP3A4:::sub::D||THBG:::ind::D
Carindacillin|ok_inv|DACA,DACB,DACC,PBPA,PBPB,MRDA,FTSI::ECOLI:inh::D|||
Procaine_benzylpenicillin|ok_vet||||
Zinc_oxide|ok||||
Zinc_sulfate|ok_inv||PPBN:::cof::D||
Sulbactam|ok|BLAT::ECOLX::6.1:C;AMPC::ENTCL::6.:C;BLA1::ECOLX::5.41:C;BLAC::STAAU:inh:5.19:DC|||
Sodium_fluoride|ok|Hydroxyapatite|A0A1C7C740:::inh::D;ENO::STRSV:inh::D;ENO::LACCB:inh::D;A0A448RWU9:::inh::D;ENOPH:::inh::D||
Ammonia_N_13|ok||NAGS:::sub::D|RHCG:::tra::D|
Tegafur_uracil|ok_inv|DPYD:::ant::D;TYSY:::ant::D;RNA;DNA|CP2A6:::sub::D;DPYD:::sub::D|S22A7:::sub::D;S29A1:::sub::D;S29A2:::sub::D;S28A1:::sub::D;S28A2:::sub::D;S28A3:::sub::D|
Vayarin|ok_inv||CP2E1:::inh::D;FADS1:::sub::D;ELOV4:::sub::D;ACOX1:::sub::D||
Antihemophilic_Factor_Recombinant_PEGylated|ok_inv|VWF:::bin::D|||VWF
Osimertinib|ok|EGFR:::inh::D|CP3A4:::duo::D;CP1A2:::ind::D|MDR1:::sub::D;ABCG2:::sub::D|
Daratumumab|ok|CD38:::abo::D|||
Kappadione|ok|THRB:::ago::D;FA7:::ago::D;FA9:::ago::D;FA10:::ago::D;PROC:::ago::D;VKGC:::ago::D;PROS:::ago::D|VKOR1:::sub::D;NCPR:::sub::D||
Iopodic_acid|ok_out|IOD3:::ant::D|||ALBU:::sub::D
Seractide_acetate|ok|ACTHR:::ago::D|||
Alatrofloxacin|ok_out||||
Technetium_Tc_99m_nofetumomab_merpentan|ok_out|EPCAM:::bin::D;CD20:::bin::D|||
Medical_air|ok_vet||||
Mersalyl|exp|PPBT:::ant::D;AQP1;MOT1:::ant::D|ITIH1:::ind::D;PCKGC:::inh::D||
Tyropanoic_acid|ok||BGLR:::sub::D||
Dextrose_unspecified_form|ok_vet||HXK1:::duo::D;HXK4:::sub_ind::D|GTR1:::sub::D;GTR2:::sub::D;GTR3:::sub::D;GLUT4:::sub::D;GTR6:::sub::D;GTR7:::sub::D;GTR8:::sub::D;GTR9:::sub::D;GTR10:::sub::D;GTR11:::sub::D;GTR12:::sub::D;SC5A1:::sub::D|
Propoxycaine|ok|CP2D6::::5.7:C;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A:::inh::D|EST1:::sub::D||
Tipiracil|ok_inv|TYPH:::inh:8.89:DC;TYPH::ECOLI::7.46:C|||S47A1:::car::DC;S22A2:::car::DC
Invert_sugar|exp||HXK4:::sub::D;PFKA::GEOSE:sub::D|GTR2:::sub::D;GTR5:::sub::D|
Pramocaine|ok|SGMR1::::7.29:C;AL1A1::::5.05:C;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A:::inh::D|||
Metrizoic_acid|ok||||
Acetrizoic_acid|out||||ALBU:::bin::D
Propiolactone|ok_out|P53::::6.6:C;DNA:::cov::D|||ALBU:::bin::D
Gastric_intrinsic_factor|ok_exp||||
Piperonyl_butoxide|ok_vet|CP3A4::::6.3:C;AL1A1::::5.:C|||
Levobetaxolol|ok_inv|ADRB1::RAT::8.3:C;ADRB1:::ant::D|CP2D6:::sub::D||
Hydroxyamphetamine|ok|TAAR1::RAT::7.3:C|||
Octasulfur|ok||||
Sulfabenzamide|ok|LMNA::::5.2:C|||
Dexpanthenol|ok||||
Rauwolfia_serpentina_root|inv|VMAT2:::inh::D|AOFA:::sub::D|SC6A2:::inh::D;Vesicle_monoamine_transporter_type_2:::inh::D|
Procaine_merethoxylline|ok||||
Propyliodone|ok||||
Polyestradiol_phosphate|ok|ESR1:::ago::D|||
Norethynodrel|ok|ANDR::RAT::5.81:C;SHBG;ANDR;ESR1|CP3A4:::sub::D||
Tannic_acid|ok||||
Trolamine_polypeptide_oleate_condensate|ok_vet||||
Indocyanine_green_acid_form|ok_inv||GLSK:::cat::D;IDHC:::cof::D|ABCBB:::sub::D;MRP2:::tra::D|
Chymotrypsin|ok_vet||||
Lapyrium|ok||||
Fluprednisolone|ok||CP3A4:::sub::D||
Sutilain|ok_out||||
Sodium_chromate_Cr_51|ok||||
Esterified_estrogens|ok||CP3A4:::sub::D||THBG:::ind::D
Meprednisone|ok_inv||CP3A5:::ind::D;CP3A4:::sub_ind::D||ALBU
Cyanocobalamin_Co_57|ok_exp||||
Norgestrel|ok|SHBG::::8.91:C;ANDR::RAT::8.37:C;GCR::::7.17:C;SC6A4::::6.23:C;LMNA::::5.55:C;ANDR:::ago::D;S5A1:::inh::D;PRGR:::bin::D|CP19A:::inh::D;CP3A4:::sub::D||
Amino_acids|inv||||
Phosphoric_acid|ok||||
Sodium_acetate|ok_inv||ACSA:::sub::D||
Technetium_Tc_99m_sulfur_colloid|ok_inv||||
Fluoride_ion_F_18|ok||||
Selenomethionine_Se_75|ok||||
Isosorbide|ok_inv|THB::::7.4:C;MCL1;B2CL1;BCL2|||
Iocetamic_acid|ok|AMPC::ECOLI::5.55:C|||
Magnesium_chloride|ok||||
Magnesium_acetate_tetrahydrate|ok|NMDA:::lig::D|||
Monopotassium_phosphate|ok_inv_vet||PPBI::BOVIN:cof:5.62:DC||
Dipotassium_phosphate|ok||||
Potassium_perchlorate|ok_inv|SC5A5:::inh::D|||ALBU:::bin::D
Xylose|ok||||
Iodide_I_123|ok||||
Protirelin|ok_inv|TRFR::MOUSE::9.31:C;TRFR::RAT::8.52:C;TRFR:::lig:8.52:DC|||
Soybean_oil|ok|PPARA:::act::D|||
Technetium_Tc_99m_polyphosphate|ok||||
Indium_In_111_pentetate|ok||||
Albumin_iodinated_I_125_serum|ok||||
Albumin_iodinated_I_131_serum|ok||||
Krypton_Kr_81m|ok||||
Safflower_oil|ok_inv||||
Technetium_Tc_99m_albumin_colloid|ok_exp||||
Sodium_phosphate_monobasic|ok|||NPT2C:::sub::D;NPT2B:::sub::D;NPT2A:::sub::D;S20A2:::sub::D;S20A1:::sub::D|
Insulin_beef|ok||CP1A2:::ind::D||
Sodium_carbonate|ok|CAH9:::inh::D;CAH4:::inh::D;CAH2:::inh::D;CAH1:::inh::D|||
Glycerin|ok_inv|LMNA::::6.45:C;TRDMT;MUTY::ECOLI:::D;RIR2::ECOLI:::D;GLPF::ECOLI:::D;MUTL::ECOLI:::D;HISX::ECOLI:::D;PAPS1;MEXA::PSEAE:::D;ARF1;ENO::ENTHR:::D;ASSY::ECOLI:::D;TGFR2;BFR::DESDA:::D;CYC4::PSEST:::D;NAGAB;PAEP;ITPR1;ADH1B;DCTD::RHIME:::D;INO1;PA2GE;GSTP1;GUNG::RUMCH:::D;HPGDS;PPARD:::ago::D|CP2E1:::ind::D;AL1A1:::sub::D||
Sodium_sulfate|ok_vet|CAH1:::inh::D;CAH2:::inh::D|||
Indium_In_111_oxyquinoline|ok||||
Enalaprilat|ok|ACE2::RAT::9.3:C;ACE::RAT::9.02:C;ACE:::inh:8.92:DC;ACE::RABIT::8.92:C;BKRB1|||
Rubidium_Rb_82|ok_inv||||ATNG:::sub::D;AT1A1:::sub::D;AT1B1:::sub::D;AT1B2:::sub::D;AT1B3:::sub::D;AT1A4:::sub::D;AT1A2:::sub::D;AT1A3:::sub::D
Iofetamine_I_123|ok||||
Magnesium_carbonate|ok_inv|NMDA:::inh::D||TRPM6:::sub::D;S41A3:::sub::D;CNNM2:::sub::D;TRPM7:::sub::D|
Potassium_lactate|ok||||
Sodium_fluorophosphate|ok||||
Iotrolan|ok||||
Acrivastine|ok|HRH1::CAVPO::5.21:C;HRH1:::ant::D|||
Indium_In_111_chloride|ok||||
Technetium_Tc_99m_red_blood_cells|ok||||
Cetyl_alcohol|ok|LMNA::::6.45:C|||
Avobenzone|ok_inv|LMNA::::7.15:C;APEX1::::5.1:C|||
Octinoxate|ok_inv||||
Strontium_chloride_Sr_89|ok_inv||PPBN:::cof::D;PPBT:::cof::D;Adenosine_triphosphate_ATP:::cof::D|NAC1:::ind::D;CAC1I:::ind::D|
Thiosulfuric_acid|ok_inv||THTR:::sub::D||
Ferric_ammonium_citrate|ok_exp||||
Fludeoxyglucose_18F|ok_inv||HXK1:::sub::D|GLUT4:::sub::D;GTR2:::sub::D;GTR1:::sub::D;GTR3:::sub::D;GTR9:::sub::D;GTR5:::sub::D;GTR6:::sub::D;GTR7:::sub::D;GTR8:::sub::D;GTR10:::sub::D;GTR11:::sub::D;GTR12:::sub::D|
Ferumoxsil|ok_exp||||
Ferumoxides|ok||||
Urea_C_13|ok|Urease::HELPY:sub::D|||
Talc|ok||||
Simethicone|ok||||
Urea_C_14|ok|Urease::HELPY:sub::D|||
Mequinol|ok||||
Sodium_ferric_gluconate_complex|ok|FRIL:::bin::D;HBA:::bin::D;HBB:::bin::D|||
Hydroquinone|ok_inv|ACES::ELEEL::8.91:C;BLM::::8.55:C;CAH2::::7.05:C;HCD2::::6.4:C;CP3A4::::6.:C;HIF1A::::5.7:C;LMNA::::5.55:C;PGDH::::5.25:C;MEN1::::5.2:C;CAH12::::5.11:C;TAU::::5.1:C;CAH3::::5.09:C;PPO2::AGABI::5.01:C;NFKB1::::5.:C;END4::ECOLI::5.:C;TYRO:::inh::D|||ALBU
Secretin_porcine|ok||||
Secretin_human|ok|SCTR:::lig:10.1:DC|||
Ecamsule|ok||||
Octocrylene|ok_inv|ESR1;ESR2|||
Titanium_dioxide|ok|MARCO|||
Iodine_povacrylex|ok||||
Omega_3_acid_ethyl_esters|ok_inv|SRBP1:::inh::D|SOAT1:::inh::D||
Methyl_salicylate|ok_vet|LMNA::::6.1:C;TSHR::::5.4:C|||
Iobenguane_sulfate_I_123|ok_inv|||SC6A2:::sub::D|
Desoxyribonuclease|ok||||
Thonzonium|ok|LMNA::::5.15:C;VATC1:::inh::D|||
Dexchlorpheniramine_maleate|ok|HRH1:::ant::D|CP3A4:::sub::D;CP2D6:::inh::D||S22A2:::inh::D;S22A1:::inh::D
Necitumumab|ok_inv|EGFR:::ant::D|||
Sodium_glycerophosphate|ok||||
Choline_C_11|ok||||
Insulin_degludec|ok|INSR:::lig::D;IGF1R|CP1A2:::ind::D||ALBU
Olive_oil|ok||||
Omega_3_carboxylic_acids|ok_inv|DGAT2:::ant::D;HCD2:::pot::D;ECHM:::pot::D;HCDH:::pot::D;ELOV4:::pot::D;LIPL:::sti::D|CP3A4:::sub::D;CP4F2:::sub::D||PPCT:::bin::D;PEBP1:::bin::D
Ixazomib|ok_inv|PSB5::::8.52:C;NFKB2::::8.21:C;PSB1::::7.51:C;PSB2::::5.46:C|CP2C9:::sub::D;CP2CJ:::sub::D;CP2D6:::sub::D;CP2C8:::sub::D;CP2B6:::sub::D;CP1A2:::sub::D;CP3A4:::sub::D||
Levmetamfetamine|ok|TAAR1::RAT::6.63:C;TAAR1::MOUSE::6.07:C;TAAR1::MACMU::5.6:C;TAAR1::::5.48:C|PNMT:::lig::D||
Clostridium_tetani|ok||||
Corynebacterium_diphtheriae|ok_inv||||
Meningococcal_groups_A_C_Y_and_W_135_oligosaccharide_diphtheria_CRM197_conjugate_vaccine|ok||||
Rabies_virus_inactivated_antigen_B|ok||||
Haemophilus_influenzae_type_B_strain_1482_capsular_polysaccharide_tetanus_toxoid_conjugate_antigen|ok_inv||||
Rotavirus_vaccine|ok||||
Rabies_virus_inactivated_antigen_A|ok_inv||||
Neisseria_meningitidis_serogroup_B_recombinant_LP2086_A05_protein_variant_antigen|ok||||
Neisseria_meningitidis_serogroup_B_recombinant_LP2086_B01_protein_variant_antigen|ok||||
Streptococcus_pneumoniae_type_4_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok_inv||||
Streptococcus_pneumoniae_type_6b_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_9v_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_14_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_18c_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_19f_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_23f_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_1_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_3_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_5_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_6a_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok_inv||||
Streptococcus_pneumoniae_type_7f_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Streptococcus_pneumoniae_type_19a_capsular_polysaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Human_papillomavirus_type_6_L1_capsid_protein_antigen|ok_inv||||
Human_papillomavirus_type_11_L1_capsid_protein_antigen|ok||||
Human_papillomavirus_type_16_L1_capsid_protein_antigen|ok_inv||||
Human_papillomavirus_type_18_L1_capsid_protein_antigen|ok_inv||||
Human_papillomavirus_type_31_L1_capsid_protein_antigen|ok||||
Human_papillomavirus_type_33_L1_capsid_protein_antigen|ok||||
Human_papillomavirus_type_45_L1_capsid_protein_antigen|ok||||
Human_papillomavirus_type_52_L1_capsid_protein_antigen|ok||||
Human_papillomavirus_type_58_L1_capsid_protein_antigen|ok||||
Measles_virus_strain_enders_attenuated_edmonston_live_antigen|ok_inv||||
Mumps_virus_strain_B_level_jeryl_lynn_live_antigen|ok_inv||||
Rubella_virus_vaccine|ok_inv||||
Varicella_Zoster_Vaccine_Live_attenuated|ok||||
Streptococcus_pneumoniae_type_1_capsular_polysaccharide_antigen|ok||||
Streptococcus_pneumoniae_type_2_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_3_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_4_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_5_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_6b_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_7f_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_8_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_9n_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_9v_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_10a_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_11a_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_12f_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_14_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_15b_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_17f_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_18c_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_19f_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_19a_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_20_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_22f_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_23f_capsular_polysaccharide_antigen|ok_inv||||
Streptococcus_pneumoniae_type_33f_capsular_polysaccharide_antigen|ok_inv||||
Haemophilus_influenzae_type_B_capsular_polysaccharide_meningococcal_outer_membrane_protein_conjugate_antigen|ok_inv||||
Bacillus_calmette_guerin_substrain_tice_live_antigen|ok||||
Ginger|ok||||
House_dust|ok||||
Acacia_longifolia_pollen|ok||||
Fraxinus_americana_pollen|ok||||
Paspalum_notatum_pollen|ok||||
Fagus_grandifolia_pollen|ok||||
Cynodon_dactylon_pollen|ok||||
Betula_lenta_pollen|ok||||
Poa_annua_pollen|ok||||
Acer_negundo_pollen|ok||||
Bromus_inermis_pollen|ok||||
Xanthium_strumarium_pollen|ok||||
Zea_mays_pollen|ok||||
Rumex_acetosella_pollen|ok||||
Rumex_crispus_pollen|ok||||
Ulmus_americana_pollen|ok||||
Ulmus_pumila_pollen|ok||||
Corylus_americana_pollen|ok||||
Carya_ovata_pollen|ok||||
Sorghum_halepense_pollen|ok||||
Poa_pratensis_pollen|ok||||
Chenopodium_album_pollen|ok||||
Acer_saccharum_pollen|ok||||
Festuca_pratensis_pollen|ok||||
Prosopis_juliflora_pollen|ok||||
Artemisia_vulgaris_pollen|ok||||
Morus_rubra_pollen|ok||||
Quercus_agrifolia_pollen|ok||||
Quercus_virginiana_pollen|ok||||
Quercus_alba_pollen|ok||||
Avena_sativa_pollen|ok||||
Olea_europaea_pollen|ok||||
Dactylis_glomerata_pollen|ok||||
Carya_illinoinensis_pollen|ok||||
Amaranthus_retroflexus_pollen|ok||||
Plantago_lanceolata_pollen|ok||||
Populus_alba_pollen|ok||||
Ambrosia_acanthicarpa_pollen|ok||||
Ambrosia_artemisiifolia_pollen|ok||||
Ambrosia_trifida_pollen|ok||||
Ambrosia_psilostachya_pollen|ok||||
Salsola_kali_pollen|ok||||
Lolium_perenne_pollen|ok||||
Artemisia_tridentata_pollen|ok||||
Atriplex_wrightii_pollen|ok||||
Platanus_occidentalis_pollen|ok||||
Platanus_racemosa_pollen|ok||||
Phleum_pratense_pollen|ok_inv||||
Holcus_lanatus_pollen|ok||||
Juglans_nigra_pollen|ok||||
Juglans_californica_pollen|ok||||
Salix_nigra_pollen|ok||||
Felis_catus_skin|ok||||
Dermatophagoides_farinae|ok||||
Dermatophagoides_pteronyssinus|ok||||
Agrostis_gigantea_pollen|ok||||
Anthoxanthum_odoratum_pollen|ok||||
Bos_taurus_skin|ok||||
Cotton_seed|ok||||
Canis_lupus_familiaris_skin|ok||||
Equus_caballus_skin|ok||||
Ceiba_pentandra_fiber|ok||||
Mus_musculus_skin|ok||||
Orris|ok||||
Rabbit|ok_inv||||
Cavia_porcellus_skin|ok||||
Periplaneta_americana|ok||||
Blatella_germanica|ok||||
Solenopsis_invicta|ok||||
Gallus_gallus_feather|ok||||
Anas_platyrhynchos_feather|ok||||
Anser_anser_feather|ok||||
Acremonium_strictum|ok||||
Alternaria_alternata|ok||||
Aspergillus_fumigatus|ok||||
Aspergillus_niger_var_niger|ok||||
Aureobasidium_pullulans_var_pullutans|ok||||
Botrytis_cinerea|ok||||
Candida_albicans|ok||||
Chaetomium_globosum|ok||||
Cladosporium_cladosporioides|ok||||
Cladosporium_sphaerospermum|ok||||
Cochliobolus_sativus|ok||||
Epicoccum_nigrum|ok||||
Fusarium_oxysporum_vasinfectum|ok||||
Helminthosporium_solani|ok||||
Mucor_plumbeus|ok||||
Neurospora_intermedia|ok||||
Penicillium_chrysogenum_var_chrysogenum|ok||||
Phoma_exigua_var_exigua|ok||||
Rhizopus_arrhizus_var_arrhizus|ok||||
Rhodotorula_rubra|ok||||
Ustilago_maydis|ok||||
Ustilago_tritici|ok||||
Stemphylium_solani|ok||||
Trichophyton_mentagrophytes|ok||||
Saccharomyces_cerevisiae|ok||||
Aspergillus_oryzae|ok||||
Aspergillus_repens|ok||||
Aspergillus_terreus|ok||||
Acacia|ok||||
Ailanthus_altissima_pollen|ok||||
Alnus_incana_subsp_rugosa_pollen|ok||||
Medicago_sativa_pollen|ok||||
Fraxinus_velutina_pollen|ok||||
Populus_tremuloides_pollen|ok||||
Morella_cerifera_pollen|ok||||
Betula_nigra_pollen|ok||||
Amaranthus_palmeri_pollen|ok||||
Juniperus_ashei_pollen|ok||||
Juniperus_virginiana_pollen|ok||||
Xanthium_strumarium_var_canadense_pollen|ok||||
Populus_deltoides_pollen|ok||||
Populus_fremontii_pollen|ok||||
Populus_deltoides_subsp_monilifera_pollen|ok||||
Cupressus_arizonica_pollen|ok||||
Taxodium_distichum_pollen|ok||||
Eupatorium_capillifolium_pollen|ok||||
Ulmus_crassifolia_pollen|ok||||
Eucalyptus_globulus_pollen|ok||||
Solidago_canadensis_pollen|ok||||
Celtis_occidentalis_pollen|ok||||
Juniperus_californica_pollen|ok||||
Robinia_pseudoacacia_pollen|ok||||
Acer_rubrum_pollen|ok||||
Melaleuca_quinquenervia_pollen|ok||||
Chenopodium_ambrosioides_pollen|ok||||
Morus_alba_pollen|ok||||
Quercus_rubra_pollen|ok||||
Syagrus_romanzoffiana_pollen|ok||||
Schinus_molle_pollen|ok||||
Amaranthus_spinosus_pollen|ok||||
Casuarina_equisetifolia_pollen|ok||||
Pinus_strobus_pollen|ok||||
Pinus_echinata_pollen|ok||||
Ligustrum_vulgare_pollen|ok||||
Elymus_repens_pollen|ok||||
Ambrosia_tenuifolia_pollen|ok||||
Ambrosia_bidentata_pollen|ok||||
Artemisia_frigida_pollen|ok||||
Distichlis_spicata_pollen|ok||||
Liquidambar_styraciflua_pollen|ok||||
Juglans_regia_pollen|ok||||
Amaranthus_tuberculatus_pollen|ok||||
Triticum_aestivum_pollen|ok||||
Felis_catus_hair|ok||||
Almond|ok||||
Apple|ok||||
Apricot|ok||||
Asparagus|ok||||
Avocado|ok||||
Banana|ok||||
Barley|ok||||
String_bean|ok||||
Beef|ok||||
Brazil_nut|ok||||
Broccoli|ok||||
Buckwheat|ok||||
Cabbage|ok||||
Cantaloupe|ok||||
Carrot|ok||||
Casein|ok||||
Celery|ok||||
Cherry|ok||||
Chicken|ok||||
Cinnamon|ok||||
Coconut|ok||||
Coffee_bean|ok||||
Red_king_crab|ok||||
Cucumber|ok||||
Egg_white|ok||||
Egg|ok||||
Egg_yolk|ok||||
Flounder|ok||||
Garlic|ok_nutra||||
Grape|ok||||
Grapefruit|ok||||
Karaya_gum|ok||||
Honeydew_melon|ok||||
Lamb|ok||||
Lemon|ok_inv||||
Lettuce|ok||||
Lima_bean|ok||||
Lobster|ok||||
Goat_milk|ok||||
Cow_milk|ok||||
Cultivated_mushroom|ok||||
Mustard_seed|ok||||
Oat|ok||||
Black_olive|ok||||
Onion|ok||||
Orange|ok||||
Oyster|ok||||
Pea|ok||||
Peach|ok||||
Peanut|ok||||
Pear|ok||||
Pecan|ok||||
Green_bell_pepper|ok||||
Black_pepper|ok||||
Pineapple|ok||||
Pistachio|ok||||
Plum|ok||||
Pork|ok||||
Potato|ok||||
Rice|ok||||
Rye|ok||||
Sesame_seed|ok||||
Shrimp|ok||||
Soybean|ok||||
Spinach|ok||||
Squash|ok||||
Strawberry|ok||||
Corn|ok||||
Tomato|ok||||
Tuna|ok||||
Turkey|ok_inv||||
Vanilla|ok||||
English_walnut|ok||||
Watermelon|ok||||
Wheat|ok||||
Tea_leaf|ok_inv||||
Khuskia_oryzae|ok||||
Artemisia_annua_pollen|ok||||
Clostridium_tetani_toxoid_antigen_formaldehyde_inactivated|ok||||
Corynebacterium_diphtheriae_toxoid_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_A_virus_A_California_7_2009_X_179A_H1N1_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Switzerland_9715293_2013_NIB_88_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Brisbane_60_2008_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_181_H1N1_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_South_Australia_55_2014_IVR_175_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_antigen_propiolactone_inactivated|ok||||
Meriones_unguiculatus_skin|ok||||
Capra_hircus_skin|ok||||
Mesocricetus_auratus_skin|ok||||
Sus_scrofa_skin|ok||||
Oryctolagus_cuniculus_skin|ok||||
Rattus_norvegicus_skin|ok||||
Bombyx_mori_fiber|ok||||
Duck|ok||||
Allergenic_extract_beef_liver|ok||||
Veal|ok||||
Bluefish|ok||||
Common_carp|ok||||
Haddock|ok||||
Pacific_halibut|ok||||
Herring|ok||||
Mackerel|ok||||
Northern_pike|ok||||
Red_snapper|ok||||
Atlantic_salmon|ok||||
European_pilchard|ok||||
Scallop|ok||||
Smelt|ok||||
Swordfish|ok||||
Trout|ok||||
White_fish|ok||||
Blackberry|ok||||
Blueberry|ok||||
Sour_cherry|ok||||
Cranberry|ok_inv||||
Date|ok||||
Fig|ok||||
Wine_grape|ok||||
Lime_citrus|ok||||
Raspberry|ok||||
Tangerine|ok||||
Artichoke|ok||||
Kidney_bean|ok||||
Beet|ok||||
Kiwi_fruit|ok||||
Brussels_sprout|ok||||
Cauliflower|ok||||
Eggplant|ok||||
Lentil|ok||||
Green_olive|ok||||
Parsley|ok||||
Sweet_potato|ok||||
Raphanus_sativus|ok||||
Rhubarb|ok||||
Turnip|ok||||
Cashew|ok||||
Hazelnut|ok||||
Macadamia_nut|ok||||
Nectarine|ok||||
Mango|ok||||
Papaya|ok||||
Leek|ok||||
Okra|ok||||
Parsnip|ok||||
Chickpea|ok||||
Black_eyed_pea|ok||||
Watercress|ok||||
Arabica_coffee_bean|ok||||
Tragacanth|ok||||
Allspice|ok||||
Laurus_nobilis|ok||||
Caraway_seed|ok||||
Clove|ok||||
Dill|ok||||
Horseradish|ok||||
Licorice|ok||||
Nutmeg|ok||||
Oregano|ok||||
Paprika|ok||||
White_pepper|ok||||
Poppy_seed|ok||||
Spearmint|ok||||
Wheat_bran|ok||||
American_chestnut|ok||||
Hops|ok||||
Musca_domestica|ok||||
Ctenocephalides_canis|ok||||
Aedes_taeniorhynchus|ok||||
Ctenocephalides_felis|ok||||
Aspergillus_flavus|ok||||
Eurotium_herbariorum|ok||||
Trichothecium_roseum|ok||||
Curvularia_inaequalis|ok||||
Fusarium_compactum|ok||||
Geotrichum_candidum|ok||||
Phoma_glomerata|ok||||
Rhodotorula_mucilaginosa|ok||||
Stemphylium_sarciniforme|ok||||
Trichoderma_harzianum|ok||||
Ustilago_avenae|ok||||
Tilletia_caries|ok||||
Puccinia_graminis|ok||||
Cotton|ok||||
Flax_seed|ok||||
Tobacco_leaf|ok||||
Corcorus_capsularis_fiber|ok||||
Agave_sisalana_fiber|ok||||
Poa_compressa_pollen|ok||||
Phalaris_arundinacea_pollen|ok||||
Bouteloua_gracilis_pollen|ok||||
Urochloa_mutica_pollen|ok||||
Secale_cereale_pollen|ok||||
Leymus_condensatus_pollen|ok||||
Pascopyrum_smithii_pollen|ok||||
Acacia_baileyana_pollen|ok||||
Alnus_rubra_pollen|ok||||
Alnus_rhombifolia_pollen|ok||||
Fraxinus_latifolia_pollen|ok||||
Betula_populifolia_pollen|ok||||
Tamarix_gallica_pollen|ok||||
Juniperus_monosperma_pollen|ok||||
Juniperus_pinchotii_pollen|ok||||
Juniperus_scopulorum_pollen|ok||||
Juniperus_osteosperma_pollen|ok||||
Juniperus_occidentalis_pollen|ok||||
Tilia_americana_pollen|ok||||
Mangifera_indica_pollen|ok||||
Acer_macrophyllum_pollen|ok||||
Acer_saccharinum_pollen|ok||||
Broussonetia_papyrifera_pollen|ok||||
Quercus_velutina_pollen|ok||||
Quercus_macrocarpa_pollen|ok||||
Quercus_kelloggii_pollen|ok||||
Quercus_gambelii_pollen|ok||||
Quercus_lobata_pollen|ok||||
Quercus_nigra_pollen|ok||||
Citrus_sinensis_pollen|ok||||
Pinus_taeda_pollen|ok||||
Pinus_palustris_pollen|ok||||
Pinus_ponderosa_pollen|ok||||
Pinus_elliottii_pollen|ok||||
Pinus_virginiana_pollen|ok||||
Pinus_monticola_pollen|ok||||
Populus_nigra_pollen|ok||||
Elaeagnus_angustifolia_pollen|ok||||
Salix_lasiolepis_pollen|ok||||
Salix_discolor_pollen|ok||||
Populus_balsamifera_subsp_trichocarpa_pollen|ok||||
Taraxacum_officinale_pollen|ok||||
Atriplex_polycarpa_pollen|ok||||
Baccharis_halimifolia_pollen|ok||||
Hymenoclea_salsola_pollen|ok||||
Allenrolfea_occidentalis_pollen|ok||||
Atriplex_lentiformis_pollen|ok||||
Artemisia_douglasiana_pollen|ok||||
Artemisia_ludoviciana_pollen|ok||||
Urtica_dioica_pollen|ok||||
Iva_axillaris_pollen|ok||||
Ambrosia_deltoidea_pollen|ok||||
Sarcobatus_vermiculatus_pollen|ok||||
Atriplex_canescens_pollen|ok||||
Artemisia_absinthium_pollen|ok||||
Japanese_encephalitis_virus_strain_sa_14_14_2_antigen_formaldehyde_inactivated|ok||||
Foreskin_fibroblast_neonatal|ok|IL6:::ago::D;VGFR1:::ago::D;IL1R1:::ago::D;TGFR2:::ago::D;FGF1:::ago::D;IFNG:::ago::D;FGFR2:::ago::D;CSF2R:::ago::D;PGFRB:::ago::D;TGFB1:::ago::D;TNFA:::ago::D|||
Bovine_type_I_collagen|ok||||
Foreskin_keratinocyte_neonatal|ok|FGF1:::ago::D;EGFR:::ago::D;CSF2R:::ago::D;IL1B:::ago::D;IL6:::ago::D;IFNG:::ago::D;FGFR2:::ago::D;PGFRA:::ago::D;TGFR2:::ago::D;TGFB1:::ago::D;TNFA:::ago::D;VEGFA:::ago::D|||
Influenza_A_virus_A_California_7_2009_H1N1_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Victoria_361_2011_H3N2_recombinant_hemagglutinin_antigen|ok||||
Influenza_B_virus_B_Wisconsin_1_2010_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Texas_50_2012_H3N2_recombinant_hemagglutinin_antigen|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Switzerland_9715293_2013_H3N2_recombinant_hemagglutinin_antigen|ok||||
Influenza_B_virus_B_Phuket_3073_2013_recombinant_hemagglutinin_antigen|ok||||
Influenza_B_virus_B_Hubei_Wujiagang_158_2009_BX_39_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Christchurch_16_2010_NIB_74_H1N1_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Victoria_361_2011_IVR_165_H3N2_antigen_propiolactone_inactivated|ok||||
Neisseria_meningitidis_serogroup_b_nhba_fusion_protein_antigen|ok||||
Neisseria_meningitidis_serogroup_b_fhbp_fusion_protein_antigen|ok||||
Neisseria_meningitidis_serogroup_b_nada_protein_antigen|ok||||
Neisseria_meningitidis_serogroup_B_strain_NZ98_254_outer_membrane_vesicle|ok||||
Bordetella_pertussis_toxoid_antigen_glutaraldehyde_inactivated|ok_inv||||
Bordetella_pertussis_filamentous_hemagglutinin_antigen_formaldehyde_inactivated|ok_inv||||
Bordetella_pertussis_pertactin_antigen|ok_inv||||
Bordetella_pertussis_fimbriae_2_3_antigen|ok_inv||||
Influenza_A_virus_A_California_7_2009_X_179A_H1N1_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_A_virus_A_Switzerland_9715293_2013_NIB_88_H3N2_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_B_virus_B_Phuket_3073_2013_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_B_virus_B_Brisbane_60_2008_antigen_formaldehyde_inactivated|ok||||
Poliovirus_type_1_antigen_formaldehyde_inactivated|ok_inv||||
Poliovirus_type_2_antigen_formaldehyde_inactivated|ok_inv||||
Poliovirus_type_3_antigen_formaldehyde_inactivated|ok_inv||||
Neisseria_meningitidis_group_a_capsular_polysaccharide_diphtheria_toxoid_conjugate_antigen|ok_inv||||
Neisseria_meningitidis_group_c_capsular_polysaccharide_diphtheria_toxoid_conjugate_antigen|ok||||
Neisseria_meningitidis_group_y_capsular_polysaccharide_diphtheria_toxoid_conjugate_antigen|ok||||
Neisseria_meningitidis_group_w_135_capsular_polysaccharide_diphtheria_toxoid_conjugate_antigen|ok||||
Influenza_A_virus_A_California_7_2009_H1N1_like_antigen_formaldehyde_inactivated|ok||||
Typhoid_Vi_polysaccharide_vaccine|ok||||
Bacillus_calmette_guerin_substrain_connaught_live_antigen|ok_inv||||
Yellow_Fever_Vaccine|ok_inv||||
Fusarium_oxysporum|ok||||
Candida_tropicalis|ok||||
Mucor_racemosus|ok||||
Penicillium_camemberti|ok||||
Penicillium_expansum|ok||||
Penicillium_italicum|ok||||
Penicillium_roqueforti|ok||||
Phoma_destructiva|ok||||
Rhizopus_stolonifer|ok||||
Fraxinus_pennsylvanica_pollen|ok||||
Atriplex_confertifolia_pollen|ok||||
Passalora_fulva|ok||||
Cochliobolus_spicifer|ok||||
Myrothecium_verrucaria|ok||||
Hypomyces_perniciosus|ok||||
Neurospora_crassa|ok||||
Paecilomyces_variotii|ok||||
Microascus_brevicaulis|ok||||
Colletotrichum_coccodes|ok||||
Pleospora_herbarum|ok||||
Streptomyces_griseus|ok||||
Trichoderma_viride|ok||||
Trichophyton_schoenleinii|ok||||
Basil|ok||||
Mung_bean|ok||||
Betula_papyrifera_pollen|ok||||
Betula_occidentalis_pollen|ok||||
Betula_alleghaniensis_pollen|ok||||
Ustilago_cynodontis|ok||||
Ustilago_nuda_hordei|ok||||
Bromus_secalinus_pollen|ok||||
Beta_vulgaris_pollen|ok||||
Chenopodium_botrys_pollen|ok||||
Mycocladus_corymbiferus|ok||||
Acrothecium_robustum|ok||||
Humicola_grisea|ok||||
Microsporum_audouinii|ok||||
Microsporum_canis|ok||||
Apiospora_montagnei|ok||||
Phycomyces_blakesleeanus|ok||||
Sporotrichum_pruinosum|ok||||
Stachybotrys_chartarum|ok||||
Syncephalastrum_racemosum|ok||||
Tetracoccosporium_paxianum|ok||||
Verticillium_albo_atrum|ok||||
White_catfish|ok||||
Carob|ok||||
Sweet_cherry|ok||||
Opilio_crab|ok||||
Bos_taurus_hair|ok||||
Serinus_canaria_feather|ok||||
Melilotus_albus_pollen|ok||||
Melilotus_officinalis_pollen|ok||||
Typha_latifolia_pollen|ok||||
Atlantic_cod|ok||||
Red_currant|ok||||
Cumin|ok||||
Cladosporium_herbarum|ok||||
Acheta_domesticus|ok||||
Canis_lupus_familiaris_hair|ok||||
Odocoileus_virginianus_hair|ok||||
Grain_mill_dust|ok||||
Epidermophyton_floccosum|ok||||
Ambrosia_dumosa_pollen|ok||||
Ambrosia_confertiflora_pollen|ok||||
Sporisorium_cruentum|ok||||
Goose|ok||||
Concord_grape|ok||||
Capra_hircus_hair|ok||||
Cavia_porcellus_hair|ok||||
Arrhenatherum_elatius_pollen|ok||||
Equus_caballus_hair|ok||||
Sus_scrofa_hair|ok||||
Carya_cordiformis_pollen|ok||||
Carya_glabra_pollen|ok||||
Millet_seed|ok||||
Mustard_greens|ok||||
Quercus_muehlenbergii_pollen|ok||||
Quercus_palustris_pollen|ok||||
Quercus_stellata_pollen|ok||||
Quercus_garryana_pollen|ok||||
Red_bell_pepper|ok||||
Perch|ok||||
Pumpkin|ok||||
Melopsittacus_undulatus_feather|ok||||
Pinus_contorta_pollen|ok||||
Pinus_sylvestris_pollen|ok||||
Pinus_rigida_pollen|ok||||
Capsicum|ok||||
Oryctolagus_cuniculus_hair|ok||||
Sequoia_sempervirens_pollen|ok||||
Rumex_obtusifolius_pollen|ok||||
Rumex_altissimus_pollen|ok||||
Rumex_salicifolius_var_mexicanus_pollen|ok||||
Sitotroga_cerealella|ok||||
English_sole|ok||||
Safflower|ok||||
Sugarcane|ok||||
Sunflower_seed|ok||||
Platanus_hybrida_pollen|ok||||
Artemisia_californica_pollen|ok||||
Helianthus_annuus_pollen|ok||||
Carpinus_caroliniana_pollen|ok||||
Picea_pungens_pollen|ok||||
Starch_tapioca|ok||||
Larix_occidentalis_pollen|ok||||
Trichophyton_rubrum|ok||||
Salix_lucida_ssp_lasiandra_pollen|ok||||
Juniperus_virginiana|ok||||
Venison|ok||||
Black_walnut|ok||||
Artemisia_dracunculus_pollen|ok||||
Pinus_banksiana_pollen|ok||||
Pinus_resinosa_pollen|ok||||
Pinus_nigra_pollen|ok||||
Pinus_thunbergii_pollen|ok||||
Carya_tomentosa_pollen|ok||||
Iva_annua_pollen|ok||||
Bassia_scoparia_pollen|ok||||
Cyclachaena_xanthifolia_pollen|ok||||
Amaranthus_retroflexus_whole|ok||||
Cephalosporium_roseum|ok||||
Cochliobolus_lunatus|ok||||
Haematonectria_haematococca|ok||||
Chrysonilia_sitophila|ok||||
Pleospora_betae|ok||||
Puccinia_striiformis_var_striiformis|ok||||
Pleospora_tarda|ok||||
Acacia_pollen|ok||||
Bassia_hyssopifolia_pollen|ok||||
Brassica_rapa_pollen|ok||||
Callistemon_citrinus_pollen|ok||||
Dicoria_canescens_pollen|ok||||
Krascheninnikovia_lanata_pollen|ok||||
Ambrosia_ambrosioides_pollen|ok||||
Ambrosia_chamissonis_pollen|ok||||
Koeleria_macrantha_pollen|ok||||
Phoenix_dactylifera_pollen|ok||||
Quercus_dumosa_pollen|ok||||
Suaeda_moquinii_pollen|ok||||
Tilia_cordata_pollen|ok||||
Apis_mellifera_venom|ok||||
Vespula_maculifrons_venom_protein|ok||||
Dolichovespula_arenaria_venom_protein|ok||||
Dolichovespula_maculata_venom_protein|ok||||
Polistes_fuscatus_venom_protein|ok||||
Hordeum_vulgare_pollen|ok||||
Agrostis_stolonifera_pollen|ok||||
Phalaris_minor_pollen|ok||||
Lolium_perenne_subsp_multiflorum_pollen|ok||||
Sorghum_bicolor_subsp_bicolor_pollen|ok||||
Sorghum_bicolor_subsp_drummondii_pollen|ok||||
Amphiachyris_dracunculoides_pollen|ok||||
Iva_angustifolia_pollen|ok||||
Neurospora_sitophila|ok||||
Trichophyton_tonsurans|ok||||
Mycogone_nigra|ok||||
Absidia_capillata|ok||||
Thermomyces_lanuginosus|ok||||
Trichosporon_cutaneum|ok||||
Tanacetum_cinerariifolium_flower|ok||||
Largemouth_bass|ok||||
Cocoa|ok||||
Blue_crab|ok||||
Barley_malt|ok||||
Radish|ok||||
Sage|ok||||
Thyme|ok||||
Peppermint|ok||||
Ulmus_rubra_pollen|ok||||
Pseudotsuga_menziesii_pollen|ok||||
Carya_laciniosa_pollen|ok||||
Maclura_pomifera_pollen|ok||||
Hepatitis_A_Vaccine|ok||||
Haemophilus_influenzae_type_B_strain_20752_capsular_polysaccharide_tetanus_toxoid_conjugate_antigen|ok_inv||||
Bordetella_pertussis_toxoid_antigen_formaldehyde_glutaraldehyde_inactivated|ok||||
Bordetella_pertussis_pertactin_antigen_formaldehyde_inactivated|ok||||
Human_papillomavirus_type_16_L1_capsid_protein_residues_2_471_antigen|ok_inv||||
Human_papillomavirus_type_18_l1_capsid_protein_residues_2_472_antigen|ok_inv||||
Influenza_A_virus_A_Christchurch_16_2010_NIB_74XP_H1N1_antigen_formaldehyde_inactivated|ok||||
Autologous_cultured_chondrocytes|ok_inv||||
Influenza_A_virus_A_Brisbane_10_2010_H1N1_antigen_MDCK_cell_derived_propiolactone_inactivated|ok_inv||||
Influenza_A_virus_A_Texas_50_2012_X_223A_H3N2_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_South_Australia_55_2014_H3N2_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Utah_9_2014_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Anthrax_vaccine|ok||||
Betula_pendula_pollen|ok||||
Ulmus_parvifolia_pollen|ok||||
Parkinsonia_florida_pollen|ok||||
Cytisus_scoparius_flowering_top|ok||||
Poultry|ok||||
Quahog_unspecified|ok||||
Cod_unspecified|ok||||
Crab_leg|ok||||
Salmon_unspecified|ok||||
Yeast|ok||||
Canis_lupus_familiaris_dander|ok||||
Cavia_porcellus_dander|ok||||
Bos_taurus_dander|ok||||
Equus_caballus_dander|ok||||
Aspergillus_nidulans|ok||||
Penicillium_digitatum|ok||||
Clonostachys_rosea_f_rosea|ok||||
Dendryphiella_vinosa|ok||||
Solenopsis_richteri|ok||||
Polistes_annularis_venom_protein|ok||||
Polistes_exclamans_venom_protein|ok||||
Polistes_metricus_venom_protein|ok||||
Vespula_germanica_venom_protein|ok||||
Vespula_pensylvanica_venom_protein|ok||||
Vespula_squamosa_venom_protein|ok||||
Vespula_vulgaris_venom_protein|ok||||
Influenza_A_virus_A_Bolivia_559_2013_H1N1_live_attenuated_antigen|ok_inv||||
Influenza_A_virus_A_Switzerland_9715293_2013_H3N2_live_attenuated_antigen|ok||||
Influenza_B_virus_B_Phuket_3073_2013_live_attenuated_antigen|ok||||
Influenza_B_virus_B_Brisbane_60_2008_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Brisbane_59_2007_H1N1_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Uruguay_716_2007_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Brisbane_60_2008_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_181_H1N1_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Victoria_210_2009_X_187_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Victoria_210_2009_X_187_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Brisbane_60_2008_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_X_223_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_BX_51B_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Switzerland_9715293_2013_NIB_88_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_H1N1_like_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Typhoid_Vaccine_Live|ok||||
Azficel_T|ok_inv||||
Human_cord_blood_hematopoietic_progenitor_cell|ok||||
Stannous_chloride|ok||||
Mineral_oil|ok_vet||||
Petrolatum|ok_inv||||
Carboxymethylcellulose|ok_inv|GTR1:::bin::D|||
Polyvinyl_alcohol|ok||||
Povidone|ok||||
Octisalate|ok_inv||||
Polysorbate_80|ok||||
Homosalate|ok_inv|PRGR:::ant::D;ANDR:::ant::D;ESR1|||
Pancrelipase_amylase|ok|Dietary_starch:::cli::D|||
Pancrelipase_protease|ok|Dietary_protein:::cli::D|||
Selenic_acid|ok||||
Phenyl_salicylate|ok|PGH2:::ant::D;PGH1:::ant::D|||
Hydrogen_fluoride|ok_inv||||
Cetylpyridinium|ok||||
Dimethicone|ok||||
Hypromellose|ok|EPCAM|||
Polyethylene_glycol_400|ok|ENPP1;HTAI2|CP4AB:::sub::D;ADHX:::sub::D;ST1A1:::sub::D||
Trolamine_salicylate|ok|PGH1:::inh::D;PGH2:::inh::D|||
Silver_nitrate|ok_inv||||
Aluminum_chloride|ok_inv|DHE3:::inh::D|||
Coal_tar|ok||||
Resorcinol|ok|LMNA::::6.:C;PGH1::SHEEP::5.44:C;CAH5B::::5.15:C;CAH12::::5.12:C;CAH2::::5.11:C;CAH5A::::5.06:C;CP3A4::::5.:C;PERT|||
Cocoa_butter|ok||||
Pyrethrum_extract|ok|NR1I2|||
Shark_liver_oil|ok||||
Docusate|ok||||
Potassium_nitrate|ok|KCNH2:::ago::D|Pentaerythritol_tetranitrate_reductase::ENTCL:sub::D|MUC1:::sub::D|
Hydrogen_peroxide|ok_vet||PPBN:::inh::D;CATA:::sub::D;GPX1:::sub::D||
Stannous_fluoride|ok||||
Calcium_Citrate|ok_inv|CASR:::ago::D;CALR:::lig::D;CIB1:::lig::D;PDCD6:::ago::D;SORCN:::lig::D;CHP1:::ago::D;SPRC:::lig::D;CALX:::lig::D;FBN2:::lig::D;S100B:::lig::D;CASQ2:::lig::D;RGN:::lig::D;PEF1:::lig::D;S10A6:::lig::D;TCTP:::lig::D;CIB2:::lig::D;S10AD:::lig::D;CASQ1:::lig::D;NUCB1:::lig::D;NUCB2:::lig::D;CALM1:::ago::D;FBN3:::lig::D;GRAN:::lig::D;CAPS1:::ago::D;CALM2:::ago::D;CALM3:::ago::D;S10AG:::lig::D;CALB2:::lig::D;CAYP1:::lig::D;CAPS2:::ago::D;CALR3:::lig::D;NRX1A:::ago::D;NCS1:::lig::D||TRPV6:::sub::D;NAC1:::sub::D;TRPV5:::sub::D;RYR1:::sub::D;RYR2:::sub::D;PK2L1:::sub::D;RYR3:::sub::D;PK1L3:::sub::D;CTSR1:::sub::D;CAC1C:::sub::D;CAC1A:::sub::D;CAC1G:::sub::D;CAC1E:::sub::D|CALB1:::sub::D;S100G:::sub::D;ALBU:::sub::D
Vitamin_D|ok_nutra_vet|VDR;VTDB|CP2R1:::sub::D;CP27B:::sub::D;CP3A4:::sub::D||
Desirudin|ok||CBPA1:::sub::D||
Meradimate|ok||||
Plantago_seed|ok_inv||||
Potassium_bicarbonate|ok|Hydrogen_ions::UNK:neu::D||S12A2:::sub::D;S12A1:::sub::D|
Allantoin|ok||||THBG:::sub::D
N_acetyltyrosine|ok||||
Sulfur_hexafluoride|ok||||
Benzalkonium|ok_inv||||
Aluminum_sesquichlorohydrate|ok||||
Magnesium_citrate|ok||||
Lanolin|ok|Skin_epithelial_cells:::coating::D|||
Castor_oil|ok_inv_nutra_vet|PE2R3:::ago::D;PE2R4:::ago::D|||
Eucalyptus_oil|ok||||
Ensulizole|ok||||
Aluminum_zirconium_trichlorohydrex_gly|ok_exp||||
Undecylenic_acid|ok_inv||||
Ammonia|ok||GLSL:::sub::D;GLNA:::sub::D;CPSM:::sub::D||
Sodium_iodide|ok||||
Turpentine|ok_exp|MK01|||
Chloroxylenol|ok|5HT2B::::5.93:C;AOFA::::5.74:C|||
Hypochlorite|ok||||
Racepinephrine|ok|ADA1A:::ago::D;ADA1B:::ago::D;ADA2A:::ago::D;ADA2B:::ago::D;ADA2C:::ago::D;ADRB1:::ago::D;ADRB2:::ago::D;ADA1D:::ant::D;ADRB3:::ago::D|||
Benzethonium|ok|LMNA::::6.7:C;RORG::MOUSE::5.4:C;CP2D6::::5.1:C;HIF1A::::5.:C|||
Calcium_gluconate|ok_vet||||
Selenious_acid|ok_inv||GPX1:::act::D;TRXR1:::sub::D|SEPP1:::tra::D|
Ammonium_molybdate|ok||||
Carbamide_peroxide|ok||||
Opium|ok_ill|OPRD:::ago::D;OPRK:::ago::D;OPRM:::ago::D|CP2D6:::sub::D;CP3A4:::sub::D||ALBU:::bin::D;B2MG:::bin::D
Capsicum_oleoresin|ok|TRPV1:::ago::D|||
Silicon_dioxide|ok|MARCO|||
Omega_3_fatty_acids|ok_nutra|PPARG:::lig::D;PPARA:::act::D;SRBP1:::inh::D|PGH2:::sub::D;LOX5:::sub::D||
Cupric_oxide|ok||||ALBU:::bin::D;CERU:::bin::D
Selenium|ok_inv_vet||SCLY:::sub::D;GSHR:::sub::D;TRXR1:::sub::D||
Chromium|ok|CYB5:::sub::D|||TRFE:::bin::D
Molybdenum|ok||||
Chromium_Cr_51|ok||||
Manganese_gluconate|ok||||
Selenomethionine|ok_inv||||
Cresol|ok||||
Oxyquinoline|ok_vet|AMPX::VIBPR::6.8:C;RORG::MOUSE::6.2:C;LEF::BACAN::6.:C;MAP2::::5.9:C|||
Aluminum_zirconium_pentachlorohydrate|ok||||
Butamben|ok_out|CP1A2::::6.5:C;LMNA::::5.15:C;CP2CJ::::5.:C;CP3A4::::5.:C;TRPV4:::inh::D;TRPA1:::inh::D;KCNJ1,KCJ10,KCJ11,KCJ12,KCJ14,KCJ15,KCNJ8:::ant::D;CCG1,CCG2,CCG3,CCG4,CCG5,CCG6,CCG7,CCG8,CA2D1,CA2D2,CA2D3,CA2D4,CAC1C,CAC1D,CAC1F,CAC1S,CACB1,CACB2,CACB3,CACB4,CAC1B,CAC1A,CAC1E,CAC1G,CAC1H,CAC1I:::inh::D|CHLE:::sub::D||ALBU:::sub::D;A1AG1:::sub::D
Aluminum_zirconium_tetrachlorohydrex_gly|ok||||
Barium_sulfate|ok||||
Sodium_hydroxide|ok||||
Trichloroacetate|ok||||
Potassium_hydroxide|ok||||
Zinc_citrate|ok||||
Triclocarban|ok|HYES::::7.89:C;HYEP::::6.92:C;EPHB::MYCTO::6.66:C;HYEP::MOUSE::6.44:C;NLRP3::::6.09:C;MEN1::::5.5:C;NPC1::::5.25:C;FABI::STAAR:ant::D|CP1B1:::ind::D;CP1A1:::ind::D||
Pyrantel|ok_vet|GPR35;ACM1:::duo::D|CP4AB:::sub::D||
Anthralin|ok|HEPS::::6.64:C;CYSP::TRYCR::6.1:C;MEN1::::6.1:C;TRYP::PIG::5.9:C;LMBL1::::5.85:C;LOX15::::5.5:C;LOX5::::5.15:C;TAU::::5.1:C;K1C12:::ant::D;JIP1:::ago::D;K22E:::ant::D|||
Pectin|ok_inv_vet||||
Sodium_sulfide|ok||||
Phenyltoloxamine|ok|DRD1::::6.46:C;DRD5::::6.38:C;DRD2::::5.56:C;DRD4::::5.56:C;HRH1::MOUSE:ANT::D|||
Polyethylene_glycol_300|ok||||
Bicisate|ok_inv||||
Rosin|ok||||
Antithrombin_Alfa|ok_inv|THRB:::inh::D;FA10:::inh::D|||
Calcium_threonate|ok||||
Ferrous_asparto_glycinate|ok||||
Ferric_sulfate|ok||||
Sesame_oil|ok_inv_nutra||||
Zinc_picolinate|ok_inv||||
Zeaxanthin|ok_inv||||
Polysorbate_20|ok||||
Exametazime|ok||||
Tetrofosmin|ok||||
Homatropine|ok|ACM5:::ant::D;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D|EST1:::sub::D||
Rose_bengal|ok_inv||LYSC:::lig::D||ALBU:::bin::D;TRFL:::bin::D;TRFE:::bin::D
Light_green_SF_yellowish|ok_exp||||
Oftasceine|ok||||
Sulisobenzone|ok|LMNA::::7.65:C;TAU::::5.25:C;Skin_epithelial_cells:::protector::D|||
Pentoxyverine|ok_inv|SGMR1::RAT::7.96:C;SGMR1:::ago:7.71:DC;PCP::::7.49:C;ACM1::::7.12:C;ACM2::::6.78:C;TSHR::::6.5:C;SC6A3::RAT::5.51:C;CP3A4::::5.4:C;CP2D6::::5.:C;OPRM:::ant::D;OPRK:::ago::D;SCN1A,SCNAA,SCNBA,SCN2A,SCN3A,SCN4A,SCN5A,SCN7A,SCN8A,SCN9A:::inh::D;KCNH2:::inh::D|||
Magnesium_glycinate|ok||||
Pantethine|ok_inv||||
Cobamamide|ok||||
Papain|ok|TLR4:::act::D|||
Ferrous_cysteine_glycinate|ok||||
Peppermint_oil|ok_inv||CP1A2:::inh::D;CP3A4:::inh::D||
Aluminum_zirconium_octachlorohydrex_gly|ok|Sweat_ducts:::ant::D|||
Menthyl_salicylate|ok|Blood_vessels:::ant::D;PGH1:::ant::D;PGH2:::ant::D|||
N_alkyl_ethylbenzyl_dimethyl_ammonium_C12_C14|ok||||
Panthenol|ok||||
Alcloxa|ok||||
Bemotrizinol|ok||||
Amiloxate|ok||||
Aluminum_chlorohydrex_propylene_glycol|ok||||
Iron_protein_succinylate|ok_inv||||
Ferrous_bisglycinate|ok||||
Arbutin|ok|TYRO:::inh::D|||ALBU
Tea_tree_oil|ok||||
Enzacamene|ok|PRGR:::ant::D;ANDR:::ant::D;ESR2;ESR1|||
Dioxybenzone|ok|SHBG:::bin::D|||FETA::RAT:bin::D
Benzoin_resin|ok||||
Peg_100_stearate|ok||||
Ethylhexyl_methoxycrylene|ok_exp||||
Methylcellulose|ok||||
Magnesium_Aluminum_Silicate|ok||||
Lycopene|ok_inv||||
Saccharide_isomerate|ok||||
Thonzylamine|ok|HRH1:::ant::D;ACM1:::ant::D;ACM2:::ant::D;ACM3:::ant::D;ACM4:::ant::D;ACM5:::ant::D|||
Trypsin|ok_vet||||
Borage_oil|ok_inv||||
Aluminum_sulfate|ok||||
Gelatin|ok_vet||||
Ethyl_macadamiate|ok||||
Cyclomethicone_5|ok||||
Copper_gluconate|ok_inv||||
Zinc_gluconate|ok_vet||||
Tocopherol|ok_inv|Free_radicals:::bin::D|CP4F2:::sub::D;CP3A4:::sub::D|TTPA:::sub::D;S14L4:::sub::D;S14L2:::sub::D;S14L3:::sub::D;APOBR:::tra::D;SCRB1:::tra::D;MDR1:::tra::D|VLDLR:::bin::D;LDLR:::bin::D
Poloxamer_407|ok_inv||||
Xanthan_gum|ok||||
Hexylresorcinol|ok|PPO2::AGABI::6.25:C;TYRO:::inh:6.25:DC;CP3A4::::5.9:C;RORG::MOUSE::5.6:C;LOX5::::5.55:C;AMPC::ECOLI::5.5:C;TAU::::5.3:C;FRIL::HORSE::5.:C;TGM2:::inh::D;TOP1:::inh::D|||
Chromium_picolinate|ok||||
Levomefolic_acid|ok_inv|SO1A3::RAT::5.92:C|METH:::cof::D|S19A1:::sub::D;PCFT:::sub::D|
Fluoride_ion|ok||||
Diacetyl_benzoyl_lathyrol|ok||||
Atractylodes_japonica_root|ok||||
Bisoctrizole|ok||||
Polydatin|ok||||
Calcium_glycerophosphate|ok||||
Sea_salt|ok||||
Protocatechualdehyde|ok|KDM4E::::5.35:C|||
Diethylamino_hydroxybenzoyl_hexyl_benzoate|ok||||
Atractylodes_japonica_root_oil|ok||||
Polysilicone_15|ok||||
Methyl_undecenoyl_leucinate|ok||||
Dihydroergocornine|ok|5HT1A:::duo::D;ADRB1:::duo::D;ADA1A:::duo::D|CP3A4:::sub::D||
Dihydro_alpha_ergocryptine|ok|DRD2:::ago::D;DRD1:::pag::D;DRD3:::pag::D|CP3A4:::sub::D||
Epicriptine|ok|DRD1:::ago::D|||
Pine_needle_oil_pinus_mugo|ok_exp||||
Aluminum_zirconium_pentachlorohydrex_gly|ok||||
DL_Methylephedrine|ok|ADRB1:::ago::D;ADA2A:::ago::D;ADA1A:::ago::D;ADRB1:::ago::D|||
Brilliant_green_cation|ok_vet|HS90A::::6.12:C;TLR9::::5.82:C|||
Diethyltoluamide|ok||||
DL_dimyristoylphosphatidylcholine|ok||||
DL_dimyristoylphosphatidylglycerol|ok||||
Ethyl_ferulate|ok_exp||||
Colloidal_oatmeal|ok_nutra||||
Rice_bran_oil|ok||||
Coccidioides_immitis_spherule|ok|HLAA:::bin::D;DRA:::bin::D;HLAA;HLAB|||
Trichophyton_verrucosum|ok||||
Thioredoxin|ok||||
Vanillyl_butyl_ether|ok||||
Thrombin|ok_inv|PAR1;PAR4;FA11:::act::D;F13A:::act::D;F13B:::act::D;FIBA:::act::D;FIBB:::act::D;FIBG:::act::D;FA5:::act::D;FA8:::act::D|||
Curcuma_aromatica_root_oil|ok||||
Hydrogenated_soybean_oil|ok||||
Phenoxyethanol|ok||||
Bentonite|ok||||
Prothrombin|ok|FIBA:::cli::D;FIBB:::cli::D;F13A:::ago::D;CBPB2:::ago::D|FA10:::sub::D||
Protein_C|ok||||
Methscopolamine|ok|ACM1::::10.02:C;ACM3::::9.87:C;ACM4::::9.85:C;ACM2::::9.75:C;ACM5::::9.68:C;ACM2:W422A:::9.36:C;ACM2:Y177Q:::9.14:C;ACM2:Y104A:::7.98:C|||
Glycol_salicylate|ok|PGH2:::ant::D;PGH1:::ant::D|||
Boric_acid|ok|LMNA::::7.35:C;TSHR::::5.8:C|||
Dipyrithione|ok|LMNA::::6.95:C;RORG::MOUSE::6.45:C;FFP::BACIU::6.15:C;HD::::5.3:C;PGH2;NOS2:::ant::D|||
Tetradecyl_hydrogen_sulfate_ester|ok|EPCR:::ant::D|||
C11_12_isoparaffin|ok||||
Factor_IX_Complex_Human|ok_inv||||
1_Palmitoyl_2_oleoyl_sn_glycero_3_phospho_rac_1_glycerol|ok_exp||||
Sinapultide|ok|Lung_epithelial_cells:::ago::D|||
Poloxamer_188|ok_inv||||
Kinetin|ok|CHIT::YEAST::5.49:C;TSHR::::5.3:C;CP1A2::::5.1:C|||
Clove_oil|ok_nutra|VCAM1:::ant::D;CXL10;CO1A1;CSF2R|||
Ubiquinol|ok_inv||||
Ichthammol|ok||||
Aluminum_oxide|ok||||
Silanol|ok||||
Rubidium|ok_inv||||
Calcium_Phosphate|ok|CASR:::ago::D;CALR:::lig::D;CIB1:::lig::D;PDCD6:::ago::D;SORCN:::lig::D;CHP1:::ago::D;SPRC:::lig::D;CALX:::lig::D;FBN2:::lig::D;S100B:::lig::D;CASQ2:::lig::D;RGN:::lig::D;PEF1:::lig::D;S10A6:::lig::D;TCTP:::lig::D;CIB2:::lig::D;S10AD:::lig::D;CASQ1:::lig::D;NUCB1:::lig::D;NUCB2:::lig::D;CALM1:::ago::D;FBN3:::lig::D;GRAN:::lig::D;CAPS1:::ago::D;CALM2:::ago::D;CALM3:::ago::D;S10AG:::lig::D;CALB2:::lig::D;CAYP1:::lig::D;CAPS2:::ago::D;CALR3:::lig::D;NRX1A:::ago::D;NCS1:::lig::D||S20A1:::sub::D;S20A2:::sub::D;NPT2A:::sub::D;NPT2B:::sub::D;NPT2C:::sub::D;TRPV6:::sub::D;NAC1:::sub::D;TRPV5:::sub::D;RYR1:::sub::D;RYR2:::sub::D;PK2L1:::sub::D;RYR3:::sub::D;PK1L3:::sub::D;CTSR1:::sub::D;CAC1C:::sub::D;CAC1A:::sub::D;CAC1G:::sub::D;CAC1E:::sub::D|CALB1:::sub::D;S100G:::sub::D;ALBU:::sub::D
Cetyl_ethylhexanoate|ok||||
Ascorbyl_phosphate|ok||||
Propolis_wax|ok||||
Polyquaternium_10_400_cps_at_2|ok||||
Linseed_oil|ok_inv||||
Guaiacol|ok|P53::::7.9:C;LEF::BACAN::6.:C;CAH2::::5.53:C;TSHR::::5.3:C;AMPC::ECOLI::5.25:C;ALBU|||
Lactobacillus_plantarum|ok_inv||||
Selexipag|ok|PI2R:::ago::D|CP3A4:::sub::D;CP2C8:::sub::D;EST1:::sub::D|MDR1:::sub::D;SO1B3:::sub::D;SO1B1:::sub::D|
Alectinib|ok_inv|ALK:::inh:8.72:DC;RET::::8.32:C;ALK:L1196M::inh:7.82:DC;VGFR2::::5.85:C||ABCG2:::inh::D|MDR1:::inh::D
Pidotimod|exp||||
Sennosides|ok|Reverse_transcriptase_RNaseH::9HIV1:inh::D;AQP3:::inh::D|||
Roquinimex|inv||||
Cefroxadine|out|PBPB::ECOLI:inh::D|BLAC::STAAU:sub::D||
Chlorophetanol|exp||||
Alfaxalone|vet|GBRP::RAT::6.52:C;GBRB2::::5.7:C;CP3A4::::5.3:C;AGAL::::5.2:C|||
Chlorobutanol|ok_inv_vet|KCNH2|||
Chloroform|ok_vet||||
Dichlorophen|exp_vet||||
Fenbendazole|vet||||
Moxidectin|ok_inv_vet|Glutamate_gated_chloride_channel::ONCVO:bin::D;GABA::ONCVO:bin::D;ABC_transporters::ONCVO:bin::D|CP3A4:::sub::D;Q14097:::sub::D|MDR1:::sub::D;ABCG2:::sub::D|
Oleandomycin|vet||CP3A4:::inh::D||
Metrifonate|vet||||
Virginiamycin|vet||||
Nalorphine|exp_vet||||
2_mercaptobenzothiazole|ok_exp_vet|PERT:::inh::D|||
Dihydrostreptomycin|inv_vet||||
Masitinib|inv_vet|ABL1::::8.68:C;ABL1:Q252H:::8.34:C;KIT:V559D-V654A:::8.33:C;KIT:V559D:::8.24:C;CSF1R::::8.12:C;KIT:L576P:::8.1:C;ABL1:F317I:::8.1:C;KIT::::8.09:C;PGFRB::::8.08:C;DDR1::::8.06:C;ABL1:F317L:::8.:C;ABL1:H396P:::7.96:C;KIT:A829P:::7.92:C;ABL1:Y253F:::7.6:C;PGFRA::::7.6:C;DDR2::::7.59:C;LCK::::7.51:C;LYN::::7.21:C;FRK::::7.06:C;ABL2::::6.96:C;ABL1:M351T:::6.85:C;FYN::::6.85:C;ABL1:E255K:::6.85:C;BLK::::6.82:C;YES::::6.24:C;FGR::::6.19:C;HCK::::6.16:C;PIM3::::6.14:C;M3K20::::6.11:C;EGFR::::6.1:C;SRC::::6.05:C;ERBB2::::5.92:C;KIT:D816V:::5.89:C;PIM1::::5.89:C;KIT:D816H:::5.82:C;RIOK2::::5.77:C;EPHA8::::5.74:C;BRAF:V600E:::5.74:C;EPHA3::::5.6:C;EGFR:L861Q:::5.33:C|||
Lesinurad|ok_inv|S22AC:::inh:5.17:DC;S22AB:::inh::D|CP3A4:::ind::D;CP2C9:::sub::D||
Aminacrine|exp|CHLE::::10.57:C;CLAT::RAT::9.82:C;CHLE::HORSE::8.92:C;ACES::ELEEL::8.7:C;ACES::::8.5:C;ACES::TETCF::8.09:C;A4::::7.91:C;ACES::MOUSE::7.74:C;ACES::BOVIN::7.57:C;AOFA::RAT::7.4:C;ACHE::::7.36:C;ACES::RAT::7.34:C;HNMT::RAT::6.96:C;ACM2::MOUSE::6.66:C;CP2D6::::6.52:C;CP1A2::::6.3:C;SC6A2::::6.29:C;S22A2::::6.17:C;S47A1::::5.96:C;ADA1A::RAT::5.95:C;ACM1::MOUSE::5.7:C;ACM2::RAT::5.68:C;NMDZ1::::5.31:C;ACM2::::5.24:C;ACM1::RAT::5.23:C;ACM2::PIG::5.2:C;SC6A4::RAT::5.12:C|||
Sebelipase_alfa|ok_inv||||
Ixekizumab|ok_inv|IL17:::abo::D|||
Padimate_O|ok|LMNA::::6.35:C;LEF::BACAN::5.3:C|||
Human_Thrombin|ok|FA5:::act::D;FA8:::act::D;FA11:::act::D;F13A:::act::D;F13B:::act::D;FIBA:::act::D;FIBB:::act::D;FIBG:::act::D|||
Thrombin_alfa|ok|FA11:::act::D;FA8:::act::D;FA5:::act::D;F13A:::act::D;F13B:::act::D;FIBA:::act::D;FIBB:::act::D;FIBG:::act::D|||
Aluminum_chlorohydrate|ok||||
Elbasvir|ok|Nonstructural_protein_5A::9HEPC:inh::D|CP343:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D|MDR1:::sub::D|
Grazoprevir|ok|Genome_polyprotein::9HEPC:ant::D|CP3A4:::sub::D|SO1B3:::sub::D;SO1B1:::sub::D;MDR1:::sub::D|A1AG1:::sub::D;ALBU:::sub::D
Ferric_oxide|exp||||
Indigotindisulfonic_acid|ok|TAU::::5.05:C;ADA1A,ADA1B,ADA1D,ADA2A,ADA2B,ADA2C:::ago::D;AHR|||
Hard_fat|ok||||
Light_Mineral_Oil|ok||||
Ravulizumab|ok_inv|CO5:::inh::D|||
Venetoclax|ok_inv|BCL2:::inh:10.44:DC;B2CL1::::7.32:C|CP3A4:::inh::D|SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|
Thiocolchicoside|exp|GABAR:::ant::D;GLRA1:::ant::D;TNF11:::ant::D|||
Cetalkonium|ok||||
Pipradrol|ok|DRD1:::ago::D|||
Drometrizole_trisiloxane|ok||||
Asunaprevir|ok_out|POLG::HCVBK:inh::D|CP2D6:::inh::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP2B6:::sub::D;CP2A6:::sub::D;CP3A5:::sub_ind::D;CP3A4:::sub_ind::D|MDR1:::inh::D;SO2B1:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D|
Etafedrine|ok|ADRB2:::ago::D|||
Carbon_monoxide|ok_inv|MYG:::deoxi::D;Alveolar_cells:::diffuse::D|||
Neon|ok_inv||||
Thimerosal|ok|METH:::ant::D;XCT:::ant::D;ATNG:::ant::D|GSHR:::ind::D;GPX1:::lig::D;SODM:::ind::D|ITPR1|ALBU
Bilastine|ok_inv|HRH1:::ant::D||SO2B1:::inh::D;SO1A2:::sub::D;ABCB5:::inh::D|
Domiphen|ok_exp||||
Atezolizumab|ok_inv|PD1L1:::abo::D|||
Levoleucovorin|ok_inv|GLYA::SHIFL:::D;DYR::ECOLI:::D|||
Human_Rho_D_immune_globulin|ok_inv|Rhesus_blood_group_D_antigen:::abo::D|||
Antithrombin_III_human|ok|ANT3:::ago::D|||
Starch_corn|ok_nutra||||
Beeswax|ok||||
Tuberculin_Purified_Protein_Derivative|ok|TLR2:::lig::D|||
Hydroxyethyl_cellulose|ok||||
Human_rabies_virus_immune_globulin|ok|GLYCO::RABVP:abo::D|||
Tetanus_Immune_Globulin|ok|TETX::CLOTE:abo::D|||
Myrrh|ok|NR1H4:::ant::D;NR1I2:::pag::D;PPARA:::ago::D|CP3A4:::ind::D||
Susoctocog_alfa|ok_inv|VWF:::bin::D|||
Efmoroctocog_alfa|ok_inv|VWF:::bin::D|||
Eftrenonacog_alfa|ok_inv||||
Normethadone|ok_ill||||
Oxilofrine|ok||||
Lifitegrast|ok|ICAM1::::8.53:C;ITAL:::ant:8.05:DC|CP2C9:::inh:5.52:DC|SO2B1:::sub::D;SO1A2:::sub::D|
Velpatasvir|ok_inv|Nonstructural_protein_5A::9HEPC:inh::D|CP2B6:::sub::D;CP2C8:::sub::D;CP3A4:::sub::D|MDR1:::inh::D;ABCG2:::inh::D;SO1B1:::inh_tra::D;SO1B3:::inh_tra::D;SO2B1:::inh_tra::D|
Rupatadine|ok|HRH1:::ant:8.41:DC;PTAFR:::ant:5.43:DC|CP2D6:::sub::D;CP2CJ:::sub::D;CP2C9:::sub::D;CP3A4:::sub::D||
Pirarubicin|inv||||
Aclarubicin|inv|5HT2B::::6.15:C;MMP2::::5.:C|||
Zorubicin|exp||||
Gestrinone|ok|SHBG:::ant:8.11:DC;ESR1:::duo::D;GNRHR:::ant::D;ANDR:::ant::D;GCR:::ant::D;PRGR:::duo::D|CP3A4:::sub::D||
Human_Varicella_Zoster_Immune_Globulin|ok||||
Dehydrocholic_acid|ok_inv|LMNA::::6.15:C|||
Epoetin_delta|ok_out||||
Perflenapent|inv_out||||
Tasonermin|ok|TNR1A:::ago::D;TNR1B:::ago::D|||
Hepatitis_B_Vaccine_Recombinant|ok_out||||
Laropiprant|ok_out|PD2R::::10.52:C;TA2R::::8.53:C;PE2R2::::6.87:C;PD2R2::::6.13:C;PE2R3::::6.05:C;PE2R1::::5.94:C;PI2R::::5.18:C;PF2R::::5.:C|||
Temoporfin|ok_inv||||
Eptotermin_Alfa|ok_out||||
Opicapone|ok_inv|COMT:::ant:9.:DC;COMT::MOUSE::8.82:C;COMT::RAT::8.82:C|CP2C8:::inh::D;CP2CJ:::ind::D||
Isavuconazole|ok_inv|CP51::CANGA:inh::D;KCNH2:::inh::D;CAC1C:::inh::D;KCNJ6:::inh::D;KCNJ9:::inh::D;KCJ11:::inh::D;KCNA5:::inh::D;KCND3:::inh::D;KCNQ1:::inh::D;SCN5A:::inh::D|CP3A4:::duo::D;CP3A5:::inh::D;CP2C8:::duo::D;CP2C9:::duo::D;CP2CJ:::inh::D;CP2D6:::inh::D;CP2B6:::ind::D;UD19:::inh::D;UD18:::inh::D|MDR1:::inh::D;ABCG2:::inh::D;S22A2:::inh::D|
Colestilan_chloride|ok_out||||
Tocofersolan|ok|MDR1:::ant::D|CP4F2:::sub::D;CP3A4:::sub::D|TTPA:::sub::D;SCRB1:::sub::D;NPCL1:::sub::D;ABCG5:::sub::D;ABCG8:::sub::D;ABCA1:::sub::D;S14L4:::sub::D;S14L2:::sub::D;S14L3:::sub::D;APOBR:::sub::D|
Nomegestrol|ok||CP3A4:::sub::D||
Delamanid|ok_inv||CP3A4:::sub::D;DDN::MYCTU:sub::D||A1AG1:::sub::D;ALBU:::sub::D
Artenimol|exp_inv|ACTG:::lig::D;AL7A1:::lig::D;ANXA2:::lig::D;ATPA:::lig::D;ATP5L:::lig::D;ATPO:::lig::D;ICAL:::lig::D;TCPG:::lig::D;COF1:::lig::D;CLIC1:::lig::D;CSRP1:::lig::D;DPYL2:::lig::D;DESP:::lig::D;EF1A1:::lig::D;ENOA:::lig::D;FLNA:::lig::D;FTO:::lig::D;G6PD:::lig::D;G3PT:::lig::D;G6PI:::lig::D;ROA2:::lig::D;HNRPD:::lig::D;HNRPK:::lig::D;HP1B3:::lig::D;HSPB1:::lig::D;IQGA1:::lig::D;FUBP2:::lig::D;LDHA:::lig::D;LDHB:::lig::D;LEG1:::lig::D;MAP4:::lig::D;MDHC:::lig::D;PSA:::lig::D;PROF1:::lig::D;PGK1:::lig::D;KPYM:::lig::D;PPIA:::lig::D;PRDX1:::lig::D;RL10:::lig::D;RL14:::lig::D;RL18:::lig::D;RL23A:::lig::D;RL35:::lig::D;RL4:::lig::D;RS13:::lig::D;RS17:::lig::D;RS18:::lig::D;RS19:::lig::D;RS28:::lig::D;RS5:::lig::D;RS6:::lig::D;RS8:::lig::D;RS9:::lig::D;SF01:::lig::D;SFPQ:::lig::D;SMD2:::lig::D;SRP14:::lig::D;SRSF4:::lig::D;TAGL:::lig::D;TAGL2:::lig::D;TPIS:::lig::D;TPM1:::lig::D;TBA1A:::lig::D;VIME:::lig::D;ZYX:::lig::D;HSP7C:::lig::D;TBB6:::lig::D;TBB4A:::lig::D;TBB5:::lig::D;ALDOA:::lig::D;G3P:::lig::D;CYC:::lig::D;PGAM1:::lig::D;MYH9:::lig::D;PDIA1:::lig::D;DDX5:::lig::D;GLYM:::lig::D;DX39B:::lig::D;NPM:::lig::D;TCTP::PLAF7:lig::D;P_type_Ca2_transporting_ATPase::PLAFA:ant::D;OAT::PLAF7:lig::D;EF1A::PLAFK:lig::D;MDR::PLAFF:lig::D;Elongation_factor_2::PLAF7:lig::D;ACT1::PLAFX:lig::D;Glyceraldehyde_3_phosphate_dehydrogenase::PLAF7:lig::D;ALF::PLAFA:lig::D;Cell_division_cycle_protein_48_homologue_putative::PLAF7:lig::D;Heat_shock_protein_90::PLAF7:lig::D;Eukaryotic_initiation_factor_4A::PLAF7:lig::D;Pyruvate_kinase::PLAF7:lig::D;LDH::PLAFD:lig::D;Protein_disulfide_isomerase::PLAF7:lig::D;Thioredoxin_related_protein_putative::PLAF7:lig::D;Spermidine_synthase::PLAF7:lig::D;Probable_ATP_dependent_6_phosphofructokinase::PLAF7:lig::D;Glutamate_dehydrogenase::PLAF7:lig::D;Endoplasmin_homolog_putative::PLAF7:lig::D;HGXR::PLAFG:lig::D;ENO::PLAF7:lig::D;40S_ribosomal_protein_S3::PLAF7:lig::D;Non::PLAF7:lig::D;TBA::PLAFK:lig::D;KNOB::PLAFA:lig::D;S_adenosylmethionine_synthase::PLAF7:lig::D;V_type_H_translocating_pyrophosphatase_putative::PLAF7:lig::D;60S_ribosomal_protein_L4::PLAF7:lig::D;Phosphoethanolamine_N_methyltransferase::PLAF7:lig::D;RS3A::PLAF7:lig::D;Conserved_Plasmodium_membrane_protein::PLAF7:lig::D;60S_ribosomal_protein_L3::PLAF7:lig::D;High_molecular_weight_rhoptry_protein_2::PLAF7:lig::D;Serine_repeat_antigen_5::PLAFA:lig::D;40S_ribosomal_protein_S19::PLAF7:lig::D;GBP::PLAF7:lig::D;ATC::PLAFK:lig::D;VATA::PLAF7:lig::D;60S_ribosomal_protein_L2::PLAF7:lig::D;Acyl_CoA_synthetase::PLAF7:lig::D;Plasmepsin_IV::PLAF7:lig::D;PLM1::PLAF7:lig::D;CRT::PLAFA:lig::D;14::PLAF7:lig::D;Isoleucine_tRNA_ligase_putative::PLAF7:lig::D;Plasmodium_exported_protein::PLAF7:lig::D;TBB::PLAF7:lig::D;60S_ribosomal_protein_L27::PLAF7:lig::D;Sec62_putative::PLAF7:lig::D;Autophagy_related_protein_18_putative::PLAF7:lig::D;Mature_parasite_infected_erythrocyte_surface_antigen::PLAF7:lig::D;Importin_7_putative::PLAF7:lig::D;Importin_subunit_alpha::PLAF7:lig::D;Peptidyl_prolyl_cis_trans_isomerase::PLAF7:lig::D;DnaJ_protein_putative::PLAF7:lig::D;MSP1::PLAFD:lig::D;Glutamate_tRNA_ligase::PLAF7:lig::D;TCPH::PLAF7:lig::D;PLM2::PLAFA:lig::D;Chaperone_putative::PLAF7:lig::D;Rhoptry_neck_protein_3::PLAF7:lig::D;40S_ribosomal_protein_S5_putative::PLAF7:lig::D;Skeleton_binding_protein_1::PLAF7:lig::D;Purine_nucleotide_phosphorylase_putative::PLAF7:lig::D;SAHH::PLAF7:lig::D;Adenosine_deaminase::PLAF7:lig::D;Methionine_tRNA_ligase::PLAF7:lig::D;Carbamoyl_phosphate_synthetase::PLAF7:lig::D;Aspartate_carbamoyltransferase::PLAF7:lig::D;Signal_recognition_particle_receptor_beta_subunit::PLAF7:lig::D;Parasite_infected_erythrocyte_surface_protein::PLAF7:lig::D;Coatomer_alpha_subunit_putative::PLAF7:lig::D;HXK::PLAFA:lig::D;Proteasome_subunit_alpha_type::PLAF7:lig::D;Haloacid_dehalogenase_like_hydrolase::PLAF7:lig::D;Insulinase_putative::PLAF7:lig::D;40S_ribosomal_protein_S21::PLAF7:lig::D;Ubiquitin_conjugating_enzyme_E2::PLAF7:lig::D;Eukaryotic_translation_initiation_factor_3_subunit_C::PLAF7:lig::D;60S_ribosomal_protein_L24_putative::PLAF7:lig::D;60S_ribosomal_protein_L23::PLAF7:lig::D;60S_ribosomal_protein_L17_putative::PLAF7:lig::D;HAP_protein::PLAF7:lig::D;Heat_shock_protein_110_putative::PLAF7:lig::D;60S_ribosomal_protein_L10_putative::PLAF7:lig::D;Lysophospholipase_putative::PLAF7:lig::D;Polyadenylate_binding_protein::PLAF7:lig::D;Ubiquitin_60S_ribosomal_protein_L40::PLAF7:lig::D;Phosphoribosylpyrophosphate_synthetase::PLAF7:lig::D;Thioredoxin_peroxidase_1::PLAF7:lig::D;Protein_transport_protein_SEC31::PLAF7:lig::D;Dipeptidyl_aminopeptidase_1::PLAF7:lig::D;RESA::PLAFF:lig::D;ATP_dependent_RNA_helicase_UAP56::PLAF7:lig::D;CDPK4::PLAF7:lig::D;RAN::PLAFA:lig::D;Nucleoside_transporter_2::PLAF7:lig::D;DRE2::PLAF7:lig::D;Glutamine_synthetase_putative::PLAF7:lig::D;60S_ribosomal_protein_L30e_putative::PLAF7:lig::D;Casein_kinase_2_alpha_subunit::PLAF7:lig::D;Threonine_tRNA_ligase::PLAF7:lig::D;cAMP_dependent_protein_kinase_regulatory_subunit::PLAF7:lig::D;Elongation_factor_1_gamma_putative::PLAF7:lig::D;Thioredoxin_like_protein::PLAF7:lig::D;60S_ribosomal_protein_L21::PLAF7:lig::D;60S_ribosomal_protein_L14_putative::PLAF7:lig::D;Inner_membrane_complex_sub_compartment_protein_3::PLAF7:lig::D;HSP40_subfamily_A_putative::PLAF7:lig::D;PDX1::PLAF7:lig::D;ALBU:::lig::D|UD19:::sub::D;UD2B7:::sub::D;CP2D6:::inh::D;CP2CJ:::inh::D||
Dibotermin_alfa|ok_inv|BMPR2:::lig::D;BMR1A:::lig::D|||
Amifampridine|ok_inv|AMPC::ECOLI::6.15:C;KCNA1:::inh::D|ARY2:::sub::D;ARY1:::sub::D||
Vinflunine|ok_inv|TBB5:::inh::D|CP3A4:::sub::D|MDR1:::sub::D;ABCB5:::sub::D|A1AG1,A1AG2:::sub::D;ALBU:::sub::D
Pitolisant|ok_inv|HRH3::CAVPO::9.8:C;HRH3:::ant:9.8:DC;HRH3::RAT::7.77:C;HRH1::::5.94:C;KCNH2:::inh::D|CP2B6:::ind::D;CP1A2:::ind::D;CP2D6:::inh::D;CP3A4:::sub_ind::D|S22A1:::inh::D|
Recombinant_Cholera_Toxin_B_Subunit|ok||||
Tafamidis|ok_inv|TTHY:::chap:8.03:DC|||
Bremelanotide|ok_inv|MC4R:::ago:9.7:DC;MSHR:::ago:8.19:DC;MC5R:::ago:7.77:DC;MC3R:::ago:7.28:DC;ACTHR:::ago::D|||
Rebamipide|inv||||
Latanoprostene_bunod|ok_inv|PF2R:::ago::D||SO2B1:::sub::D|
Curcumin|ok_exp_inv|LEF::BACAN::7.1:C;CISD1::::7.:C;PTGES::::6.7:C;NPSR1::::6.5:C;AOFA::::6.15:C;A4::::5.82:C;LMNA::::5.75:C;PGH1::BOVIN::5.7:C;SRC::MOUSE::5.66:C;TAU::::5.52:C;HD::::5.45:C;MEN1::::5.4:C;HCD2::::5.4:C;HIF1A::::5.2:C;EP300::::5.19:C;FRIL::HORSE::5.15:C;TLR9::::5.08:C;EGFR::::5.06:C;AL1A1::::5.05:C;ABHD5::::5.04:C;TSHR::::5.:C;CBR1;MRP5:::inh::D;VDR;PPARG|GSTM1:::inh::D;GSTA1:::inh::D;CP2D6:::inh::D;CP1A2:::inh::D;CP2B6:::inh::D;CP3A4:::inh::D;CP2C9:::inh::D;GSTP1:::inh::DC|MDR1:::inh::D|
Treosulfan|inv||||
Naldemedine|ok_inv|OPRM:::ant::D;OPRD:::ant::D;OPRK:::ant::D|CP3A4:::sub::D;UD13:::sub::D|ABCB5:::sub::D|
Voclosporin|inv|CANB1;CANB2|||
Racecadotril|inv||||
Ipragliflozin|inv|SC5A2::::8.13:C|||
Tropisetron|ok_inv|5HT3A:::ant:10.6:DC;5HT3A::RAT::9.22:C;5HT3B::MOUSE::8.42:C;5HT1A::::8.28:C;ACHA7::::8.16:C;ACHA7::MOUSE::8.16:C;ACHA7::RAT::8.:C;5HT3A::CAVPO::7.52:C;5HT4R::CAVPO::7.27:C;5HT4R::RAT::7.2:C;5HT4R::::6.7:C;SC6A4::::6.59:C;CP3A4::::6.3:C;ACHB4::::5.74:C;ACM5::::5.61:C;ACM1::RAT::5.35:C|||
Acalabrutinib|ok_inv|BTK:::inh::D|CP3A4:::inh::D;CP3A5:::inh::D;CP3A4:::sub::D||ALBU:::bin::D;A1AG1:::bin::D
Iomeprol|ok_inv||||
Tezacaftor|ok_inv|CFTR:::act::D|CP3A4:::sub::D;CP3A5:::sub::D|MDR1:::inh::D|
Durvalumab|ok_inv|PD1L1:::bin::D;CD80:::bin::D|||
Epacadostat|inv||||
Encorafenib|ok_inv|BRAF:V600E::inh:9.52:DC;BRAF:::inh:9.52:DC;MK14::::5.66:C;CCND1:::inh::D|CP2D6:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D||
Ribociclib|ok_inv|CDK4:::ant::D;CDK6:::ant::D|CP3A4:::inh::D||
Lasmiditan|ok_inv|5HT1F:::ago::D|CP2D6:::inh::D|MDR1:::inh::D;ABCG2:::inh::D;S22A1:::inh::D;S47A1:::inh::D;S47A2:::inh::D|
Galactose|ok_inv||||
Icotinib|exp_inv|EGFR:::ant:8.7:DC|CP3A5:::sub_ind::D;CP1A2:::sub::D;CP3A4:::sub::D||
Rilmenidine|ok_inv|NISCH::RAT::7.95:C;ADA2C::::7.9:C;ADA2A::::7.44:DC;ADA2B::::7.37:C;NISCH::::7.23:C;CP2D6::::6.4:C;ADA1A::::5.22:C;CP3A4::::5.1:C;CP2C9::::5.:C|||
Ebastine|ok_inv|HRH1::::8.48:C;5HT2A::::7.59:C;ADA2C::::7.4:C;DRD3::::7.38:C;HRH1::CAVPO::7.35:C;5HT1A::::7.33:C;DRD2::::7.21:C;SC6A3::::7.11:C;KCNH2::::7.07:C;ACM1::::6.99:C;ACM4::::6.94:C;5HT2C::::6.91:C;ACM3::::6.86:C;ADA1A::::6.74:C;5HT2B::::6.7:C;ADA1B::RAT::6.63:C;ACM5::::6.61:C;ACM2::::6.55:C;ADA2A::::6.51:C;ADA2B::::6.47:C;DRD4::::6.34:C;SC6A2::::6.34:C;EGFR::::6.25:C;DRD1::::6.22:C;SC6A4::::6.19:C;NK2R::::6.19:C;FYN::::6.09:C;ADA1D::::6.06:C;5HT6R::::5.99:C;ERBB2::::5.98:C;ADA1A::RAT::5.98:C;5HT1B::RAT::5.85:C;MDR1::::5.82:C;AA3R::::5.74:C;ADRB3::::5.72:C;HRH2::::5.54:C;MTOR::::5.33:C;LMNA::::5.2:C;ACES::::5.13:C|CP3A4:::sub::D||
Benfotiamine|ok_exp||||
Clobetasol|ok_exp_inv||CP3A5:::ind::D;CP3A4:::sub_ind::D||
Rifamycin|ok_inv|RPOB::ECOLI:bin::D;RPOA::ECOLI:bin::D;RPOC::ECOLI:bin::D|CP3A4:::duo::D;CP2CJ:::duo::D;CP2B6:::duo::D;CP2C8:::duo::D;CP2C9:::duo::D;CP1A2:::inh::D|SO1A2:::inh::D;SO1B1:::inh::D;SO1B3:::inh::D;SO2A1:::inh::D;SO2B1:::inh::D;S47A1:::inh::D;MDR1:::inh::D|ALBU:::sub::D
Istradefylline|ok_inv|AA2AR::RAT::8.7:C;AA2AR:::ant:8.66:DC;AA1R::RAT::6.82:C;AA1R:::ant:6.08:DC;AA2BR::::5.74:C;AA3R::::5.35:C|CP2D6:::sub::D;CP2CI:::sub::D;CP2C9:::sub::D;CP2C8:::sub::D;CP2B6:::sub::D;CP1A2:::sub::D;CP3A4,CP343,CP3A5,CP3A7:::inh::D;CP3A5:::sub::D;CP3A4:::sub::D;CP1A1:::sub::D|S47A2:::inh::D;S47A1:::inh::D;PO2F2:::inh::D;S22A6:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Talazoparib|ok_inv|PARP1:::inh:9.24:DC;PARP2:::inh:9.07:DC||ABCG2:::sub::D;MDR1:::sub::D|
Tenapanor|ok_inv|SL9A3:::inh:8.3:DC;SL9A3::RAT::8.03:C|CP3A5:::sub::D;CP3A4:::sub::D||
Sarilumab|ok_inv|IL6RA:::aab::D;FCGR1;FCG2A;FCG2B;FCG3A;FCG3B|ALAT1:::ind::D;ALAT2:::ind::D;Aspartate_aminotransferase:::ind::D;CP3A4:::duo::D||
Zytron|ok_inv||||
Talinolol|inv||CP2D6:::sub::D||
Pazufloxacin|inv|STRP::STRP1::5.21:C|CP1A2:::inh::D||
Brodalumab|ok_inv||||
Imidapril|inv|ACE::::5.:C|||
Neuropeptide_Y|ok_inv||||
Capmatinib|ok_inv|MET::::9.89:C|||
Niraparib|ok_inv|PARP1:::ant:8.7:DC;PARP2:::ant:8.68:DC;PARP4::::6.48:C;TNKS1::::6.24:C;PARP3::::5.89:C|BGLR:::sub::D;Q6LAP9:::sub::D||
Aceneuramic_acid|inv||||
Bictegravir|ok_inv|Reverse_transcriptase_RNaseH::9HIV1:ant::D;Integrase::9HIV1:ant::D|CP3A4:::sub::D;UD11:::sub::D;PO2F2:::inh::D;S47A1:::inh::D||
Tivozanib|inv|VGFR2::::9.8:C;VGFR1::::9.68:C;VGFR3::::9.62:C;PGFRA::::8.65:C;EPHB2::::7.76:C|||
Sirukumab|inv||||
Faldaprevir|inv|SOAT2::RAT::5.62:C;PP2BB::::5.05:C|||
Tilarginine|ok_inv|NOS2::::8.74:C;NOS1::RAT::7.:C;NOS3::::6.52:C;NOS1::::6.08:C;NOS2::MOUSE::5.64:C;NOS1::MOUSE::5.37:C;NOS3::BOVIN::5.15:C|||
Baricitinib|ok_inv|JAK2:::inh:9.1:DC;JAK1:::inh:9.:DC;TYK2::::8.06:C;JAK3:::inh:7.6:DC;FAK2:::inh::D|CP3A4:::sub::D|SO1B3:::inh::D;S22A2:::inh::D;S22A6:::inh::D;S47A2:::inh::D;ABCG2:::inh::D;S22A8:::inh::D|
Nifurtimox|inv||||
Esketamine|ok_inv|NMDZ1::::7.94:C;NMDZ1::RAT::6.19:C;NTRK2;BDNF:::ago::D;EF2:::inh::D;NMDE2:::ant::D;NMDA:::ant::D|CP2C9:::sub::D;CP2CJ:::sub::D;CP3A4:::sub_ind::D;CP2B6:::sub_ind::D||
Ertugliflozin|ok_inv|SC5A4::::9.06:C;SC5A2::RAT::8.94:C;SC5A1::::5.71:C;SC5A2:::ant::D|UD14:::inh::D;UD11:::inh::D;UD2B7:::sub::D;UD19:::sub::D|ABCG2:::sub::D;MDR1:::sub::D|ALBU:::bin::D
Neratinib|ok_inv|EGFR:::inh:10.1:DC;EGFR:G719C::inh:9.43:DC;EGFR:L861Q::inh:9.43:DC;M4K5::::9.19:C;EGFR:L858R::inh:9.17:DC;EGFR:G719S::inh:9.04:DC;ERBB2::::9.:C;EGFR:T790M::inh:8.82:DC;ERBB4::::8.62:C;STK24::::8.19:C;STK26::::8.13:C;M4K3::::8.11:C;ERBB3::::8.11:C;STK25::::7.92:C;STK10::::7.89:C;MP2K1::::7.85:C;M3K19::::7.8:C;MP2K2::::7.59:C;EGFR:L858R-T790M::inh:7.57:DC;MINK1::::7.54:C;M3K4::::7.41:C;STK3::::7.24:C;MP2K5::::7.2:C;SLK::::7.18:C;PAK2::::7.1:C;BLK::::7.07:C;M4K1::::7.03:C;E2AK4::::7.02:C;LCK::::6.92:C;M3K3::::6.89:C;TNIK::::6.85:C;NUAK2::::6.85:C;BTK::::6.8:C;UFO::::6.72:C;PAK1::::6.68:C;M4K2::::6.66:C;SIK1::::6.66:C;YES::::6.62:C;GAK::::6.6:C;NEK2::::6.6:C;STK4::::6.57:C;KC1E::::6.54:C;M4K4::::6.48:C;ST17A::::6.47:C;M3K12::::6.43:C;TIE1::::6.41:C;MERTK::::6.4:C;M3K2::::6.35:C;HCK::::6.31:C;FER::::6.29:C;MP2K7::::6.28:C;CSK::::6.26:C;FES::::6.23:C;CSF1R::::6.17:C;ACK1::::6.17:C;M3K13::::6.13:C;LYN::::6.09:C;KPCD1::::6.09:C;VGFR2::::6.07:C;CHK2::::6.07:C;STK33::::6.03:C;ST17B::::5.96:C;KPCD2::::5.96:C;WEE2::::5.89:C;NUAK1::::5.82:C;M3K20::::5.82:C;HIPK4::::5.82:C;MELK::::5.8:C;FGR::::5.72:C;FAK1::::5.72:C;JAK3::::5.7:C;CDK16::::5.64:C;IRAK1::::5.64:C;KPCD3::::5.62:C;NEK3::::5.62:C;MK10::::5.6:C;EPHB6::::5.55:C;INSR::::5.52:C;TIE2::::5.52:C;FLT3:D835Y:::5.51:C;SIK2::::5.48:C;MK08::::5.48:C;MET::::5.4:C;SRC::::5.39:C;WEE1::::5.39:C;KS6A2::::5.39:C;TAOK3::::5.38:C;MET:Y1235D:::5.38:C;STK35::::5.35:C;FLT3:D835H:::5.34:C;INSRR::::5.34:C;M3K10::::5.34:C;TXK::::5.32:C;FLT3:K663Q:::5.31:C;CDK7::::5.29:C;KSYK::::5.29:C;STK36::::5.28:C;FLT3::::5.27:C;M3K9::::5.27:C;MAST1::::5.26:C;KCC1D::::5.25:C;CHK1::::5.24:C;M3K11::::5.24:C;ABL1:Q252H:::5.22:C;FLT3:N841I:::5.19:C;ST32B::::5.19:C;FYN::::5.19:C;DUSTY::::5.19:C;KC1G2::::5.18:C;MET:M1250T:::5.17:C;KS6A1::::5.13:C;PAK6::::5.12:C;KC1G3::::5.11:C;FAK2::::5.1:C;RON::::5.08:C|FMO3:::sub::D;CP3A4:::sub::D|MDR1:::inh::D|A1AG1,A1AG2:::sub::D;ALBU:::sub::D
Guselkumab|ok_inv|IL23A:::inh::D|||
Indium_In_111_pentetreotide|ok_inv||||
Angiotensin_II|ok_inv|AGTR2::::10.1:C;AGTRB::RAT::10.:C;AGTR1:::ago:9.8:DC;AGTRA::RAT::9.4:C;AGTR1::BOVIN::8.24:C|||
Revefenacin|ok_inv|ACM1:::ant::D|CP2D6:::sub::D|SO1B1:::sub::D;SO1B3:::sub::D;MDR1:::sub::D;ABCG2:::sub::D|ALBU:::bin::D
Brexanolone|ok_inv|GBRA1::::7.66:C;GBRP::RAT::7.29:C;GBRA5::MOUSE::6.06:C;NPSR1::::5.5:C;MEN1::::5.1:C;GEMI::::5.:C;GABAR:::aga::D|ALDR:::sub::D||
Romosozumab|ok_inv|SOST:::inh::D|||
Alanyl_glutamine|inv||||
Prulifloxacin|inv||CP1A2:::inh::D||
Apalutamide|ok_inv|ANDR:::ant:7.46:DC;GABAR:::ant::D|CP2C9:::ind::D;CP2CJ:::ind::D;CP2C8:::sub::D;CP3A4:::sub_ind::D|S47A1:::inh::D;S47A2:::inh::D;S22A8:::inh::D;S22A2:::inh::D;SO1B1:::ind::D;ABCG2:::ind::D;MDR1:::ind::D|
Rociletinib|inv||||
Valbenazine|ok_inv|Vesicle_monoamine_transporter_type_2:::ant::D|CP2D6:::sub::D;CP3A4:::sub::D;CP3A5:::sub::D||
Deflazacort|ok_inv|GCR:::ago::D|CP3A5:::ind::D;CP3A4:::sub_ind::D||
Flomoxef|inv||||
Selinexor|ok_inv|XPO1:::inh::D|CP3A4:::sub::D|SO1B3:::inh::D|
Delafloxacin|ok_inv|PARC::ECOLI:inh::D;GYRA::ECOLI:inh::D|UD11:::sub::D;UD13:::sub::D;UDB15:::sub::D;CP2E1:::ind::D;CP2C9:::ind::D;CP3A4:::ind::D|ABCB5:::sub::D;ABCG2:::sub::D|ALBU:::sub::D
Avelumab|ok_inv|PD1L1:::ant::D|||
Lemborexant|ok_inv|OX1R:::ant::D;OX2R:::ant::D|CP3A4:::sub::D;CP3A5:::sub::D;CP2B6:::ind::D;CP3A4:::duo::D|MDR1:::sub::D|
Duvelisib|ok_inv|PK3CG:::inh:8.54:DC;PK3CD:::inh::D|CP3A4:::sub::D|ABCG2:::sub::D;MDR1:::sub::D|
Dacomitinib|ok_inv|ERBB2::::9.2:C;EGFR:::inh:8.74:DC;ERBB4::::7.13:C;LCK::::7.03:C;SRC::::6.96:C;JAK3::::5.45:C|UD11:::inh::D;CP2C9:::sub::D;CP3A4:::sub::D;CP2D6:::inh::D|S22A1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|ALBU:::bin::D
Binimetinib|ok_inv|MP2K2:::inh::D;M3K1:::inh::D;IL1B;TNFA;IL6|CP2CJ:::sub::D;CP1A2:::sub::D;UD11:::sub::D||
Glasdegib|ok_inv|SMO::MOUSE::8.3:C;SMO:::inh::D|UD19:::sub::D;CP2C8:::sub::D;CP3A4:::sub::D|S47A2:::inh::D;S47A1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|ALBU:::sub::D
Elagolix|ok_inv|GNRHR|CP3A4:::sub::D;CP2D6:::sub::D;CP2C8:::sub::D|MDR1:::sub::D;SO1B1:::sub::D|
Entrectinib|ok_inv|NTRK1:::inh:9.:DC;ALK::::9.:C;LTK::::8.8:C;NTRK3:::inh:8.8:DC;NTRK2:::inh:8.6:DC;ROS1:::inh:8.3:DC;FER::::8.3:C;FRK::::7.8:C;JAK2:::inh:7.7:DC;SRC::::7.5:C;ACK1::::7.5:DC;RET::::7.4:C;UFO::::7.4:C;CSF1R::::7.4:C;PLK4::::7.4:C;IGF1R::::7.2:C;FAK1::::7.:C;JAK1::::6.95:C;FGFR3::::6.8:C;KIT::::6.8:C;BTK::::6.8:C;SLK::::6.8:C;FLT3::::6.79:C;PTK6::::6.71:C;BLK::::6.7:C;LYN::::6.7:C;VGFR3::::6.7:C;CLK4::::6.7:C;INSR::::6.68:C;AURKA::::6.67:C;RON::::6.6:C;FGFR1::::6.6:C;AAPK1::::6.6:C;ABL1::::6.5:C;AURKB::::6.47:C;JAK3::::6.46:C;M4K2::::6.4:C;FYN::::6.4:C;VGFR2::::6.4:C;LCK::::6.3:C;KSYK::::6.2:C;KPCG::::6.2:C;M4K5::::6.2:C;VGFR1::::6.1:C;MET::::6.1:C;CLK2::::6.:C;KS6A3::::5.9:C;PKN2::::5.9:C;CDK7::::5.9:C;HIPK2::::5.8:C;KPCT::::5.8:C;STK3::::5.7:C;M4K4::::5.7:C;TBK1::::5.6:C;KCC1D::::5.6:C;DAPK3::::5.6:C;LRRK2::::5.6:C;GRK5::::5.6:C;TAOK1::::5.5:C|CP3A4:::sub::D|MDR1:::inh::D|
Ocrelizumab|ok_inv|CD20:::aab::D|||
Benznidazole|ok_inv|AMPC::ECOLI::5.25:C|||
Diacerein|ok_inv|TAU::::5.55:C;GLD1::CAEEL::5.14:C;CASP3::::5.1:C;HS90A::::5.03:C;RORG::MOUSE::5.:C;MEN1::::5.:C;CP2D6:::inh::D;CP2C9:::inh::D;CP2E1:::inh::D;CP3A4,CP343,CP3A5,CP3A7:::inh::D;CP1A2:::inh::D;LOX5:::inh::D;Arylamine_N_acetyltransferase::HELPY:inh::D;NR1H2:::inh::D;NR1H3:::inh::D|||
Avatrombopag|ok_inv|ABCG2:::inh::D;TPOR:::ago::D;S22A8:::inh::D|CP2C8:::ind::D;CP2C9:::ind::D|MDR1:::sub::D|
Thymopentin|inv||||
Vosaroxin|inv||||
Abemaciclib|ok_inv|CDK4:::inh:9.22:DC;CCND3::::8.09:C;CCND1::::8.:C;CCNT1::::7.24:C;CDK1::::6.43:C;CDK5::::6.39:C;CCNE1::::6.3:C;CCNH::::5.51:C;CDK6:::inh::D|CP2D6:::inh::D;CP2C9:::inh::D;CP2C8:::inh::D;CP2B6:::inh::D;CP1A2:::inh::D;CP3A4:::inh::D|MDR1:::inh::D;ABCG2:::inh::D;S22A2:::inh::D;S47A2:::inh::D;S47A1:::inh::D|A1AG1,A1AG2:::bin::D;ALBU:::bin::D
Fostamatinib|ok_inv|KSYK:::inh:7.77:DC;ST32A:::inh::D;ST17B:::inh::D;ST17A:::inh::D;STK16:::inh::D;STK10:::inh::D;SRMS:::inh::D;SRC:::inh::D;SNRK:::inh::D;SLK:::inh::D;SIK2:::inh::D;SIK1:::inh::D;SGK3:::inh::D;SBK3:::inh::D;SBK1:::inh::D;KS6A3:::inh::D;KS6A1:::inh::D;ROS1:::inh::D;ROCK2:::inh::D;RIPK4:::inh::D;RIPK2:::inh::D;RIPK1:::inh::D;RIOK3:::inh::D;RIOK2:::inh::D;RIOK1:::inh::D;RET:::inh::D;RAF1:::inh::D;PTK6:::inh::D;FAK2:::inh::D;FAK1:::inh::D;PRP4B:::inh::D;KGP2:::inh::D;KPCD1:::inh::D;KPCT:::inh::D;KPCI:::inh::D;KPCG:::inh::D;KPCE:::inh::D;KPCD:::inh::D;KAPCB:::inh::D;AAPK1,AAPK2,AAKB1,AAKB2,AAKG1,AAKG2,AAKG3:::inh::D;AAPK1:::inh::D;PLK4:::inh::D;PLK3:::inh::D;PLK2:::inh::D;PLK1:::inh::D;PKN2:::inh::D;PKN1:::inh::D;PMYT1:::inh::D;PI42C:::inh::D;PI42B:::inh::D;PIM3:::inh::D;PIM1:::inh::D;PK3CG:::inh::D;PK3CD:::inh::D;P3C2G:::inh::D;P3C2B:::inh::D;PI4KB:::inh::D;PHKG1:::inh::D;CDK15:::inh::D;PDPK1:::inh::D;PGFRB:::inh::D;PGFRA:::inh::D;CDK17:::inh::D;CDK16:::inh::D;PAK5:::inh::D;PAK6:::inh::D;PAK4:::inh::D;PAK3:::inh::D;PAK2:::inh::D;PAK1:::inh::D;OXSR1:::inh::D;NUAK2:::inh::D;NUAK1:::inh::D;NTRK3:::inh::D;NTRK2:::inh::D;NTRK1:::inh::D;NEK9:::inh::D;NEK5:::inh::D;NEK4:::inh::D;NEK3:::inh::D;NEK2:::inh::D;NEK11:::inh::D;NEK1:::inh::D;MYO3A:::inh::D;MYLK4:::inh::D;MYLK3:::inh::D;MYLK2:::inh::D;MYLK:::inh::D;MUSK:::inh::D;RON:::inh::D;MKNK2:::inh::D;MKNK1:::inh::D;MINK1:::inh::D;MERTK:::inh::D;MELK:::inh::D;MATK:::inh::D;MAST1:::inh::D;CLAP1:::inh::D;MARK4:::inh::D;MARK3:::inh::D;MARK2:::inh::D;MARK1:::inh::D;MAPK5:::inh::D;MK09:::inh::D;MK07:::inh::D;MK04:::inh::D;MK15:::inh::D;MK14:::inh::D;MK13:::inh::D;MK10:::inh::D;M4K5:::inh::D;M4K4:::inh::D;M4K3:::inh::D;M4K2:::inh::D;M4K1:::inh::D;M3K9:::inh::D;M3K6:::inh::D;M3K4:::inh::D;M3K3:::inh::D;M3K2:::inh::D;M3K15:::inh::D;M3K13:::inh::D;M3K12:::inh::D;M3K11:::inh::D;M3K10:::inh::D;M3K1:::inh::D;MP2K6:::inh::D;MP2K5:::inh::D;MP2K3:::inh::D;MP2K2:::inh::D;LYN:::inh::D;LTK:::inh::D;LRRK2:::inh::D;LIMK2:::inh::D;LIMK1:::inh::D;LCK:::inh::D;LATS1:::inh::D;KIT:::inh::D;SIK3:::inh::D;VGFR2:::inh::D;JAK3:::inh::D;JAK2:::inh::D;ITK:::inh::D;IRAK4:::inh::D;IRAK3:::inh::D;IRAK1:::inh::D;INSRR:::inh::D;INSR:::inh::D;IKKE:::inh::D;IKKB:::inh::D;ICK:::inh::D;HIPK3:::inh::D;HIPK2:::inh::D;HCK:::inh::D;GSK3B:::inh::D;GSK3A:::inh::D;GAK:::inh::D;FYN:::inh::D;FRK:::inh::D;MTOR:::inh::D;VGFR3:::inh::D;FLT3:::inh::D;VGFR1:::inh::D;FGR:::inh::D;FGFR3:::inh::D;FGFR2:::inh::D;FGFR1:::inh::D;FES:::inh::D;FER:::inh::D;ERN1:::inh::D;ERBB4:::inh::D;ERBB2:::inh::D;EPHB6:::inh::D;EPHB4:::inh::D;EPHB2:::inh::D;EPHB1:::inh::D;EPHA8:::inh::D;EPHA7:::inh::D;EPHA6:::inh::D;EPHA5:::inh::D;EPHA4:::inh::D;EPHA3:::inh::D;EPHA2:::inh::D;EPHA1:::inh::D;E2AK4:::inh::D;E2AK2:::inh::D;E2AK1:::inh::D;EGFR:::inh::D;DYR1B:::inh::D;DYR1A:::inh::D;DDR2:::inh::D;DDR1:::inh::D;DCLK3:::inh::D;DCLK2:::inh::D;DCLK1:::inh::D;DAPK3:::inh::D;DAPK2:::inh::D;DAPK1:::inh::D;CSK22:::inh::D;CSK21:::inh::D;KC1A:::inh::D;CSK:::inh::D;CSF1R:::inh::D;CLK4:::inh::D;CLK3:::inh::D;CLK2:::inh::D;CLK1:::inh::D;CTRO:::inh::D;CHK2:::inh::D;CHK1:::inh::D;CDKL2:::inh::D;CDKL1:::inh::D;CDK4:::inh::D;MRCKG:::inh::D;CDK1:::inh::D;CASK:::inh::D;CSKP:::inh::D;KKCC2:::inh::D;KKCC1:::inh::D;KCC2G:::inh::D;KCC2D:::inh::D;KCC2B:::inh::D;KCC2A:::inh::D;KCC1G:::inh::D;KCC1D:::inh::D;KCC1A:::inh::D;BTK:::inh::D;BRAF:::inh::D;BMX:::inh::D;BMPR2:::inh::D;BMR1B:::inh::D;BMP2K:::inh::D;BLK:::inh::D;UFO:::inh::D;AURKC:::inh::D;AURKB:::inh::D;AURKA:::inh::D;ANKK1:::inh::D;ALK:::inh::D;COQ8B:::inh::D;ACV1B:::inh::D;ACVR1:::inh::D;ABL2:::inh::D;AAK1:::inh::D;ZAP70:::inh::D;M3K20:::inh::D;M3K19:::inh::D;YES:::inh::D;WEE1:::inh::D;ULK3:::inh::D;ULK2:::inh::D;ULK1:::inh::D;TYRO3:::inh::D;TXK:::inh::D;TTK:::inh::D;TSSK1:::inh::D;TNI3K:::inh::D;ACK1:::inh::D;TNK1:::inh::D;TNIK:::inh::D;TLK2:::inh::D;TLK1:::inh::D;TIE1:::inh::D;TGFR2:::inh::D;TGFR1:::inh::D;TESK1:::inh::D;TIE2:::inh::D;TBK1:::inh::D;TAOK3:::inh::D;TAOK2:::inh::D;TAOK1:::inh::D;STK39:::inh::D;ST38L:::inh::D;STK38:::inh::D;STK36:::inh::D;STK35:::inh::D;STK33:::inh::D;TEC:::inh::D;STK3:::inh::D;STK24:::inh::D;KAPCA:::inh::D;STK26:::inh::D;NIM1:::inh::D;MET:::inh::D;JAK1:::inh::D;COQ8A:::inh::D;TYK2:::inh::D;KS6A6:::inh::D;PKNB::MYCTU:inh::D;CDPK1::PLAF7:inh::D;ABL1:::inh::D;CATL1:::inh::D;CATS:::inh::D;LOX5:::inh::D;PDE5A:::inh::D;UD11:::inh::D;S29A1:::inh::D;FAAH1:::inh::D;Vesicle_monoamine_transporter_type_2:::inh::D;AA3R:::ant::D|UD19:::sub::D;CP3A4:::inh::D|ABCB5:::sub::D;ABCG2:::inh::D|
Alpelisib|ok_inv|PK3CA:::inh:8.34:DC;PK3CG::::6.6:C;PK3CD::::6.54:C;PK3CB::::5.92:C;PK3CB::RAT::5.66:C|CP2CJ:::inh::D;CP2C8:::inh::D;CP2C9:::ind::D;CP3A4:::sub::D|MDR1:::inh::D;ABCG2:::sub::D|
Tecovirimat|ok_inv|F13::VAR67:inh::D|UD11:::sub::D;UD14:::sub::D||
Benralizumab|ok_inv|IL5RA:::abo::D;FCG3A:::bin::D|||
Voxilaprevir|ok_inv|Genome_polyprotein::9HEPC:inh::D|CP3A4:::sub::D;CP1A2:::sub::D;CP2C8:::sub::D|MDR1:::inh::D;ABCG2:::inh::D;SO1B1:::inh::D;SO1B3:::inh::D|
Sarecycline|ok_inv|||MDR1:::inh::D|
Letermovir|ok_inv|TRM3::HCMVM:inh::D;TRM2::HCMVM:inh::D;TRM1::HCMVM:inh::D|CP343:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::inh::D;CP2B6:::ind::D;CP2C9:::ind::D;CP2CJ:::ind::D;CP2C8:::inh::D;CP2D6:::sub::D;UD13:::sub::D;UD11:::sub::D|MRP2:::inh::D;S22A8:::inh::D;ABCBB:::inh::D;ABCG2:::inh::D;MDR1:::inh::D;SO1B3:::sub::D;SO1B1:::sub::D|
Gefarnate|inv||||
Anecortave|inv||||
Oxitropium|inv||||
Gadolinium|ok_inv||||
Telotristat_ethyl|ok_inv|TPH2:::ant::D;TPH1:::ant::D|||
Mannitol_busulfan|ok_inv||||
Vaborbactam|ok_inv|AMPC::ENTCL:inh::D;BLKPC::KLEPN:inh::D;Beta_lactamase::KLEPN:inh::D;Q939N4,Q9L5C7,Q840M4:::inh::D;Beta_lactamase::ECOLX:inh::D;BLA1::KLEPN:inh::D;BLAT::ECOLX:inh::D;Beta_lactamase::KLEPN:inh::D;Beta_lactamase::KLEPN:inh::D|||
Cinepazide|inv||||
Sultamicillin|ok_inv||||
Lorlatinib|ok_inv|ALK:F1174L::inh:9.7:DC;ALK:L1196M::inh:9.15:DC;ALK:::inh:8.89:DC;ALK:C1156Y::inh:8.8:DC;LTK::::8.57:C;FER::::8.48:C;ALK:S1206Y::inh:8.38:DC;FES::::8.22:C;ALK:L1152R::inh:8.05:DC;FAK2::::7.85:C;ALK:G1269A::inh:7.82:DC;ACK1::::7.77:C;FAK1::::7.77:C;NTRK2::::7.64:C;NTRK1::::7.62:C;NTRK3::::7.34:C;FRK::::7.28:C;ALK:G1202R::inh:7.11:DC|UD13:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP2B6:::ind::D;CP3A5:::sub::D;CP3A4,CP343,CP3A5,CP3A7:::inh::D||
Vinpocetine|inv|BLM::::6.1:C;HIF1A::::5.2:C;TAU::::5.05:C|CP3A4:::sub::D||
Gilteritinib|ok_inv|FLT3:::inh:9.39:DC;ALK:::inh:8.82:DC;ROS1::::8.72:C;RET::::8.47:C;UFO:::inh::D;5HT1A,5HT1B,5HT1D,5HT1E,5HT1F,5HT2A,5HT2B,5HT2C,5HT3A,5HT3B,5HT3C,5HT3D,5HT3E,5HT4R,5HT6R,5HT7R:::inh::D|CP3A4:::sub::D|S22A1:::inh::D;ABCG2:::inh::D;S47A1:::inh::D;MDR1:::sub::D|ALBU:::bin::D
Erdafitinib|ok_inv|FGFR1:::inh::D;FGFR2:::inh::D;FGFR3:::inh::D;FGFR4:::inh::D;RET_proto_oncogene:::sub::D;CSF1R:::sub::D;PGFRA:::sub::D;PGFRB:::sub::D;KIT:::sub::D;VGFR2:::sub::D|CP2C9:::sub::D;CP3A4:::sub::D|MDR1:::inh::D;S22A2:::inh::D|
Citicoline|ok_exp|LicC_protein::STRPN:::D|||
Dupilumab|ok_inv|IL4RA:::ant::D|||
Bucillamine|inv||||
Deutetrabenazine|ok_inv|VMAT2:::inh::D|CBR1:::sub::D;CBR3:::sub::D;CP2D6:::sub::D;CP1A2:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D||
Nimorazole|inv||||
Gepirone|inv|5HT1A::::7.89:C;5HT1A::RAT::7.5:C;DRD2::::7.24:C;ADA1B::RAT::5.62:C|||
Faropenem|inv||||
Iron_isomaltoside_1000|ok_inv||||
Landiolol|inv||CP2D6:::sub::D||
Bergapten|inv|DYR1A::RAT::5.83:C;CP2D6::::5.7:C;CP2CJ::::5.5:C;TSHR::::5.4:C;CP2C9::::5.3:C;CP3A4::::5.:C|||
Canrenone|inv||||
Polatuzumab_vedotin|ok_inv|CD79B|CP3A4:::sub::D|CD79B|
Edaravone|ok_inv|LEF::BACAN::8.8:C;KDM4E::::5.95:C;AL1A1::::5.6:C;DNAB::MYCTU::5.56:C;TAU::::5.55:C;RECA::MYCTU::5.53:C||S22A8:::sub::D;S22A6:::sub::D|
Triclabendazole|ok_inv|STRP::STRP1::5.53:C;HS90A::::5.37:C;TAU::::5.1:C;MEN1::::5.:C;Q6IX08,CYSB,CATLL,CATL1,CATL2,ENO,K7YNB3,NU3M::FASHE:inh::D|CP2B6:::inh::D;CP2C8:::inh::D;CP2A6:::inh::D;CP2D6:::inh::D;CP2CJ:::inh::D;CP1B1:::sub::D;CP1A1:::sub::D;CP3A4:::inh::D;CP2C9:::sub::D;CP1A2:::inh::D||
Tulobuterol|inv|ADRB2::BOVIN::6.89:C;ADRB2|||
Stem_bromelain|ok_inv||||
Moxaverine|inv||||
Fexinidazole|inv||||
Brigatinib|ok_inv|ALK:::inh::D;EGFR:::inh::D;ABL1:::inh::D;IGF1R:::inh::D;FLT3:::inh::D;INSR:::bin::D;MET:::inh::D;ERBB4:::inh::D;ERBB2:::inh::D|CP2C8:::sub::D;CP3A4:::sub::D;CP3A4:::ind::D|ABCB5:::inh::D;ABCG2:::inh::D;S22A1;S47A1:::inh::D;S47A2:::inh::D|
Polihexanide|ok_inv||||
Propiverine|ok_inv|ADA1A:::ant::D;CAC1C:::ant::D;ACM5;ACM4:::ant::D;ACM3:::ant::D;ACM2:::ant::D;ACM1:::ant::D|FMO3:::sub::D;FMO1:::sub::D;CP3A4:::sub::D||
Luspatercept|ok_inv||||
Nefopam|ok_inv||||
P_nitrobiphenyl|ok_exp_inv||||
Doravirine|ok_inv|Reverse_transcriptase_RNaseH::9HIV1:inh::D|CP3A5;CP3A4:::sub::D||
Dopexamine|ok_inv||||
Benzbromarone|inv_out|CP2C9:::inh:8.1:DC;S22AC::::7.66:C;LMNA::::7.35:C;AK1C1::::7.32:C;MRP1::::6.72:C;UBP2::::6.2:C;HIF1A::::6.:C;5HT2B::::5.94:C;MK14::::5.91:C;MK01::::5.71:C;DNAB::MYCTU::5.56:C;AA3R::::5.53:C;TSHR::::5.4:C;CP2J2::::5.37:C;S22A6::::5.34:C;PPARG::::5.32:C;STRP::STRP1::5.18:C|CP2CJ:::inh:5.43:DC|ABCBB:::sub::D;SO2B1:::inh::D;SO1B1:::inh::D|
Cantharidin|ok_inv|PPM1B::::6.37:C;LMNA::::5.95:C;PP1G::::5.75:C;HIF1A::::5.6:C;PTN1::::5.44:C;RORG::MOUSE::5.3:C;MK01::::5.3:C;Skin_epithelial_cells:::ves::D;AHR:::ago::D|||
Eravacycline|ok_inv|RS4::ECOLI:inh::D|AOFA:::sub::D;CP3A4:::sub::D||
Rucaparib|ok_inv|PARP1:::ant:9.09:DC;TNKS2::::7.85:C;TNKS1::::7.6:C;DYR1A::::6.3:C;PIM1::::5.9:C;CDK1::::5.6:C;KPCD2::::5.3:C;PARP3:::ant::D;PARP2:::ant::D|UD11:::inh::D;CP2C8:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D;CP343:::inh::D;CP3A7:::inh::D;CP3A5:::inh::D;CP3A4:::idw::D;CP1A2:::duo::D;CP2D6:::inh::D|S22A8:::inh::D;S22A6:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;MRP4:::inh::D;S22A1:::inh::D;S47A2:::inh::D;S47A1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|
Carisbamate|inv||||
Temocillin|ok_inv||||
Diaminopropanol_tetraacetic_acid|ok_inv||||
Betrixaban|ok_inv|FA10:::inh:9.93:DC|THRB:::inh::D|KCNH2:::inh:5.74:DC;MDR1:::sub::D|
Vestronidase_alfa|ok_inv||||
Siponimod|ok_inv|S1PR1::::9.4:DC;S1PR5:::mod:9.01:DC;S1PR4::::6.12:C;S1PR3::::5.3:C|CP2C9:::sub::D;CP3A4:::sub::D||
Velmanase_alfa|inv||||
Relebactam|ok_inv|AMPC::ENTCL:inh::D;Beta_lactamase::KLEPN:inh::D;Q939N4,Q9L5C7,Q840M4:::inh::D;BLA1::ECOLX:inh::D;BLAT::ECOLX:inh::D||S47A2:::sub::D;S47A1:::sub::D;S22AB:::sub::D;S22A8:::sub::D|
Polmacoxib|inv||||
Bromperidol|ok_inv|CP2D6::::5.4:C;CP1A2::::5.3:C;AMPC::ECOLI::5.1:C;CP3A4::::5.:C|||
Iobitridol|ok_inv||||
Gemigliptin|inv||||
Steviolbioside|ok_inv||||
Nadifloxacin|inv|LMNA::::6.15:C|||
Omadacycline|ok_inv|RS3::ECOLI:inh::D;RS7::ECOLI:inh::D;RS8::ECOLI:inh::D;RS19::ECOLI:inh::D;RS14::ECOLI:inh::D;16S_ribosomal_RNA::Gut_flora:inh::D||MDR1:::sub::D|ALBU
Ketanserin|inv|5HT2A::RAT::9.55:C;5HT2A:::ANT:9.55:DC;5HT2B::RAT::9.4:C;SGMR1::::9.:C;5HT2C::RAT::8.92:C;5HT2A::PIG::8.88:C;HRH1::CAVPO::8.85:C;HRH1::::8.7:C;AA3R::::8.57:C;DRD4::::8.46:C;ADA1B::RAT::8.09:C;5HT2C::::7.36:C;5HT2B::::6.74:C;DRD2::::6.62:C;5HT1D::::6.59:C;AL1A1::::6.45:C;DRD2::RAT::6.44:C;PGDH::::6.25:C;5HT1A::::6.1:C;5HT7R::::5.87:C;5HT1A::RAT::5.74:C;5HT1B::RAT::5.72:C;CP2CJ::::5.6:C;LMNA::::5.6:C;5HT6R::::5.55:C;CP2C9::::5.4:C;5HT1B::::5.19:C|||
Levodropropizine|inv||||
Taurolidine|ok_inv||||
Lynestrenol|ok_inv||CP3A4:::sub::D;CP2C9:::sub::D;CP2CJ:::inh::D||
Piribedil|inv|NFKB1::::6.95:C;CP2D6::::6.7:C;CP2CJ::::6.2:C;CP1A2::::5.7:C;CP3A4::::5.5:C;ACM1::RAT::5.05:C;DRD3;DRD2|||
Copanlisib|ok_inv|PK3CA:::inh:9.3:DC;PK3CD:::inh:9.15:DC;PK3CB::::8.43:C;PK3CG::::8.19:C|CP343:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub::D|S47A2:::inh::D;ABCG2:::sub::D;MDR1:::sub::D|ALBU:::sub::D
Promestriene|inv||||
Piritramide|ok_inv||||
Mogamulizumab|ok_inv|CXCR4:::ant::D|||
Fedratinib|ok_inv|GAK::::8.96:C;JAK2:::inh:8.96:DC;DAPK3::::8.92:C;FLT3:D835H::inh:8.31:DC;FLT3:D835Y::inh:8.19:DC;STK16::::8.18:C;DCLK3::::7.89:C;FLT3:::inh:7.89:DC;FLT3:K663Q::inh:7.89:DC;DAPK1::::7.8:C;JAK1:::inh:7.74:DC;M3K19::::7.72:C;FLT3:N841I::inh:7.7:DC;TYK2::::7.68:C;DAPK2::::7.54:C;FLT3:R834Q::inh:7.54:DC;BMP2K::::7.49:C;NUAK1::::7.47:C;AAK1::::7.46:C;FYN::::7.42:C;SIK1::::7.41:C;ABL1:E255K:::7.4:C;FAK1::::7.38:C;ABL1::::7.36:C;PGFRB::::7.35:C;ST17B::::7.35:C;ABL1:H396P:::7.35:C;KIT:A829P:::7.34:C;RET::::7.32:C;NUAK2::::7.31:C;ABL1:M351T:::7.3:C;ABL1:Q252H:::7.27:C;ABL1:Y253F:::7.25:C;KIT:V559D:::7.24:C;ACK1::::7.19:C;ABL1:T315I:::7.19:C;PI51A::::7.18:C;MK07::::7.18:C;RET:V804L:::7.15:C;LCK::::7.14:C;JAK3::::7.13:C;SRC::::7.12:C;ULK2::::7.1:C;RET:V804M:::7.09:C;FGR::::7.09:C;TBK1::::7.04:C;RIOK3::::7.04:C;PLK4::::7.02:C;SIK2::::7.01:C;RIOK1::::7.:C;PKNB::MYCTU::7.:C;SRPK2::::7.:C;E2AK4::::7.:C;YES::::6.92:C;IRAK3::::6.92:C;NEK6::::6.92:C;KIT:L576P:::6.92:C;CDK7::::6.92:C;CSK22::::6.92:C;KIT::::6.89:C;MYLK4::::6.89:C;CTRO::::6.85:C;KS6A4::::6.85:C;RET:M918T:::6.82:C;NEK9::::6.82:C;ACVR1::::6.82:C;NEK7::::6.8:C;KIT:D816H:::6.8:C;KIT:D816V:::6.8:C;UFO::::6.8:C;PI42B::::6.8:C;SRPK1::::6.8:C;BRD4::::6.79:C;SRPK3::::6.77:C;GRK4::::6.77:C;ABL1:F317L:::6.74:C;DCLK1::::6.72:C;FRK::::6.7:C;MK10::::6.7:C;STK33::::6.66:C;HIPK4::::6.66:C;FAK2::::6.66:C;IRAK1::::6.66:C;SNRK::::6.64:C;MK09::::6.62:C;MK08::::6.59:C;ULK1::::6.57:C;FGFR1::::6.55:C;PLK1::::6.55:C;ULK3::::6.54:C;COQ8B::::6.52:C;KCC2A::::6.52:C;MARK3::::6.52:C;EPHB6::::6.52:C;STK11::::6.51:C;PHKG1::::6.48:C;BRDT::::6.47:C;AURKC::::6.46:C;CDK17::::6.46:C;IKKE::::6.44:C;KS6A6::::6.44:C;MP2K5::::6.44:C;FGFR3::::6.44:C;IKKB::::6.44:C;TNK1::::6.44:C;MKNK2::::6.42:C;WEE1::::6.41:C;PRP4B::::6.41:C;BMR1B::::6.39:C;KS6A1::::6.38:C;TTK::::6.35:C;KCC1D::::6.34:C;FGFR2::::6.33:C;ITK::::6.31:C;AURKB::::6.31:C;LYN::::6.3:C;MK15::::6.29:C;MYLK::::6.28:C;FES::::6.28:C;KCC2G::::6.27:C;ABL1:F317I:::6.25:C;M3K2::::6.24:C;NEK5::::6.24:C;ABL2::::6.24:C;EGFR:L858R-T790M:::6.24:C;EGFR:T790M:::6.24:C;KCC2D::::6.23:C;M3K13::::6.23:C;ROS1::::6.22:C;ST17A::::6.21:C;CSF1R::::6.21:C;M3K20::::6.19:C;BLK::::6.19:C;NEK3::::6.19:C;ALK::::6.19:C;SLK::::6.17:C;TIE1::::6.15:C;MARK1::::6.15:C;EPHA1::::6.14:C;TAOK2::::6.12:C;FGFR3:G697C:::6.12:C;MUSK::::6.1:C;SBK1::::6.1:C;MERTK::::6.09:C;NTRK1::::6.08:C;IKKA::::6.08:C;HIPK1::::6.07:C;BTK::::6.07:C;INSR::::6.07:C;STK36::::6.06:C;LRRK2::::6.06:C;CDK4::::6.06:C;DCLK2::::6.06:C;CSK21::::6.04:C;LIMK1::::6.03:C;DDR2::::6.02:C;MARK4::::6.01:C;E2AK1::::6.:C;HIPK2::::6.:C;LRRK2:G2019S:::6.:C;DMPK::::6.:C;PKN1::::5.96:C;FER::::5.96:C;E2AK2::::5.96:C;TGFR2::::5.96:C;PTK6::::5.92:C;IRAK4::::5.92:C;PAK5::::5.92:C;NEK11::::5.92:C;CDPK1::PLAF7::5.92:C;ERN1::::5.92:C;BMX::::5.92:C;MK06::::5.92:C;HIPK3::::5.89:C;TLK1::::5.89:C;TAOK1::::5.89:C;TSSK1::::5.89:C;M4K1::::5.89:C;M3K3::::5.89:C;CDKL2::::5.89:C;KIT:V559D-T670I:::5.82:C;TXK::::5.82:C;EGFR::::5.82:C;KGP2::::5.8:C;STK39::::5.8:C;INSRR::::5.8:C;PHKG2::::5.8:C;KCC1A::::5.8:C;PLK3::::5.8:C;NEK4::::5.8:C;DUSTY::::5.77:C;MATK::::5.77:C;NEK2::::5.77:C;EPHB1::::5.77:C;PI4KB::::5.77:C;TNI3K::::5.74:C;KKCC1::::5.74:C;M4K3::::5.74:C;ICK::::5.72:C;TAOK3::::5.72:C;SIK3::::5.72:C;TIE2::::5.72:C;DDR1::::5.72:C;CLK4::::5.7:C;FGFR4::::5.7:C;TLK2::::5.7:C;ERBB4::::5.7:C;VGFR3::::5.7:C;KS6B1::::5.7:C;ROCK1::::5.68:C;HCK::::5.68:C;EPHB4::::5.68:C;M4K2::::5.68:C;IGF1R::::5.66:C;KS6A5::::5.66:C;ROCK2::::5.66:C;KS6A2::::5.64:C;CLK2::::5.64:C;PLK2::::5.62:C;AAPK1::::5.62:C;ACVL1::::5.62:C;SGK3::::5.6:C;CLK1::::5.6:C;CDK14::::5.59:C;MELK::::5.59:C;RIOK2::::5.59:C;GRK7::::5.59:C;PGFRA::::5.57:C;CDK18::::5.57:C;KSYK::::5.57:C;CSKP::::5.55:C;STK10::::5.54:C;SBK3::::5.54:C;BMPR2::::5.54:C;MYLK2::::5.52:C;NTRK2::::5.51:C;CDK16::::5.51:C;MARK2::::5.51:C;MP2K2::::5.51:C;M3K7::::5.51:C;M3K11::::5.51:C;PAK1::::5.51:C;TESK1::::5.49:C;KCC1G::::5.49:C;M3K9::::5.49:C;EGFR:L858R:::5.48:C;NEK1::::5.47:C;KIT:V559D-V654A:::5.46:C;MP2K3::::5.46:C;KGP1::::5.42:C;ZAP70::::5.42:C;PAK4::::5.42:C;CHK1::::5.42:C;PK3CA:H1047L:::5.41:C;EPHB2::::5.41:C;EPHA6::::5.41:C;KKCC2::::5.4:C;EPHA4::::5.4:C;M3K4::::5.39:C;PI42C::::5.39:C;ANKK1::::5.37:C;VGFR1::::5.37:C;NIM1::::5.36:C;MET:M1250T:::5.36:C;AURKA::::5.36:C;EPHA2::::5.36:C;AAPK2::::5.33:C;SRMS::::5.3:C;MP2K1::::5.29:C;VGFR2::::5.28:C;RIPK1::::5.28:C;STK38::::5.24:C;EGFR:L861Q:::5.24:C;CSK::::5.23:C;WEE2::::5.22:C;PAK2::::5.22:C;RIPK2::::5.21:C;M3K12::::5.2:C;LTK::::5.2:C;EPHA7::::5.19:C;KCC2B::::5.17:C;ACV1B::::5.17:C;PAK6::::5.16:C;M3K10::::5.16:C;COQ8A::::5.15:C;EPHA3::::5.15:C;STK25::::5.14:C;MKNK1::::5.14:C;CDKL5::::5.14:C;STK26::::5.12:C;PK3CG::::5.12:C;EPHA8::::5.11:C;LIMK2::::5.1:C;LATS2::::5.1:C;KPCE::::5.09:C;KS6A3::::5.09:C;CDK15::::5.07:C;NTRK3::::5.07:C;MET::::5.07:C;CDK9::::5.06:C;MINK1::::5.05:C;BRAF:V600E:::5.03:C;KPCD3::::5.02:C;DYR1B::::5.02:C;RIPK4::::5.01:C;MYLK3::::5.01:C;BRAF::::5.01:C;MP2K4::::5.:C|FMO3:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D|S47A2:::inh::D;S47A1:::inh::D;PO2F2:::inh::D;SO1B3:::inh::D;SO1B1:::inh::D;ABCG2:::inh::D;MDR1:::inh::D|
Mizolastine|ok_inv|HRH1::::8.57:C;KCNH2::::6.46:C|CP2D6:::inh::D||
Molgramostim|inv||||
Nitrite|ok_inv||||
Oxetacaine|ok_inv|LMNA::::7.35:C;SCN1A::::5.64:C;CP2D6::::5.5:C;HIF1A::::5.1:C;GAST:::inh::D|CP3A4:::inh:5.1:DC||
Benzodiazepine|ok_inv||CP3A4:::sub::D||
Indobufen|inv||||
Mebeverine|ok_inv||||
Pentetreotide|ok_inv||||
Sisomicin|inv||||
Ozanimod|inv||||
Plazomicin|ok_inv|RS14::ECOLI:inh::D;30S_ribosomal_protein_S11::ENTBF:inh::D||S47A1:::inh::D;S47A2:::inh::D|
Octenidine|inv||||
Evogliptin|inv|DPP4::::9.05:C|||
Somatorelin|inv||||
Urapidil|inv|LMNA::::6.3:C;CP2CJ::::5.1:C|||
Protionamide|ok_inv|LMNA::::6.1:C;PPO2::AGABI::5.35:C|||
Moxetumomab_Pasudotox|ok_inv|CD22:::bin::D;EF2:::inh::D|||
Gusperimus|inv||||
Ibalizumab|ok_inv|CD4:::ant::D;CCR5:::ant::D;CXCR4:::ant::D|||
Balugrastim|inv||||
Sulprostone|inv|RORG::MOUSE::5.6:C;MEN1::::5.:C|||
Perazine|ok_inv||||
Fenpropidin|ok_exp||||
Iodide|ok_exp|CAH5B::::7.6:C|||
Cicletanine|inv||||
Gaxilose|ok_inv||||
BCG_vaccine|inv||||
Lafutidine|inv||||
Benserazide|ok_inv|DDC:::inh::D|||
Norethandrolone|inv||||
Dinoprost|ok_inv|PF2R::::8.6:C;PF2R::MOUSE::7.9:C;SO2A1::::7.64:C;SO2A1::RAT::7.35:C;SO2A1::MOUSE::6.98:C;PE2R3::::6.96:C;PF2R::BOVIN::6.89:C;PE2R1::::6.66:C;SO2B1::RAT::6.54:C;TA2R::::5.85:C;PE2R4::::5.38:C;PD2R::::5.35:C;PD2R2:::ago::D|||
Boscalid|ok_exp||||
Trifarotene|ok_inv|RARG:::ago::D;RARB:::ago::D;RARA:::ago::D|CP2C9:::sub::D;CP3A4:::sub::D;CP2C8:::sub::D;CP2B6:::sub::D||
Cepeginterferon_alfa_2B|inv||CP1A2:::inh::D||
Perflubutane|ok_inv||||
Lefamulin|ok_inv|RL22::STRPN:bin::D|CP3A4:::sub:5.35:DC|MDR1:::sub::D|
Amithiozone|inv||||
Prednimustine|inv||||
Secnidazole|ok|MK01::::5.3:C;ATM::::5.15:C|||
Pegvaliase|ok_inv||||
Reproterol|inv||||
Melarsoprol|inv||||
Etelcalcetide|ok_inv|CASR:::ago::D|||
Benperidol|ok_inv|DRD2::::10.57:C;DRD4::::10.18:C;DRD3::::9.54:C;5HT2A::::8.92:C;HIF1A::::6.1:C;LMNA::::5.8:C;CP2D6::::5.2:C|||
Vonicog_Alfa|ok_inv|FA8:::stbz::D;CO1A1:::bin::D|ATS13:::sub::D||
Oxatomide|inv|HRH1::CAVPO::8.05:C;KPYM::::7.6:C;DRD3::::7.2:C;NR1I2::::6.4:C;CP2D6::::6.1:C;LEF::BACAN::5.9:C;MEN1::::5.5:C;ACM1::RAT::5.3:C;CP2C9::::5.1:C;HIF1A::::5.:C|||
Trofosfamide|inv||||
Factor_XIII_human|ok_inv||||
Nicoboxil|ok_inv||||
Gallopamil|inv|CAC1C::::7.77:C;LMNA::::6.25:C;MDR1::::5.49:C;SCN1A::::5.44:C|CP3A4:::sub::D||
Ozenoxacin|ok_inv|GYRA::HAEIN:inh::D;PARC::ECOLI:inh::D|||
Cafedrine|inv||||
Theodrenaline|inv||||
Opipramol|inv|SGMR1::::9.7:C;EBP::::7.89:C;ERG2::YEAST::7.77:C|||
Isoxaflutole|ok_exp_inv||||
Darolutamide|ok_inv|ANDR:::ant::D;PRGR:::ant::D|CP3A4:::sub::D;UD19|ABCG2:::inh::D;MDR1:::sub::D|ALBU:::bin::D
Lactitol|inv||||
Phloroglucinol|inv||||
Dihydralazine|ok_exp||CP1A2:::inh::D||
Pivagabine|inv||||
Methylprednisone|ok_inv||CP3A4:::sub::D||
Terizidone|ok_inv||||
Prothipendyl|inv||||
Silver|ok_inv|MTF1:::bin::D;CERU:::bin::D;ALBU:::bin::D;A2MG:::bin::D|||
Mitoguazone|inv||||
Pyronaridine|inv||||
Pexidartinib|ok_inv|CSF1R:::inh::D;KIT:::inh::D;FLT3:::inh::D;PGFRB:::inh::D|CP3A4:::duo::D;UD14:::sub::D;CP2B6:::duo::D;CP2C9:::inh::D;UD11:::inh::D|S47A1:::inh::D;S47A2:::inh::D;SO1B1:::inh::D;SO1B3:::inh::D;SO2B1:::inh::D|ALBU:::bin::D;A1AG1:::bin::D
Silicon|ok_inv||||
Cortivazol|inv|GCR|CP3A4:::ind::D;CP3A5:::ind::D||
Enfortumab_vedotin|ok_inv|NECT4:::bin::D|CP3A4:::sub::D|MDR1:::sub::D|
Tiapride|inv|LMNA::::8.15:C;ACM1::RAT::6.45:C;DRD3:::inh:6.41:DC;DRD2:::inh:6.39:DC;ADA2A,ADA2B,ADA2C:::ant:6.11,,:DC;ADA2A::::6.11:C;TSHR::::5.2:C;CP2D6::::5.1:C;ADA1A,ADA1B,ADA1D:::ant::D;5HT1A,5HT1B,5HT1D,5HT1E,5HT1F,5HT2A,5HT2B,5HT2C,5HT3A,5HT3B,5HT3C,5HT3D,5HT3E,5HT4R,5HT6R,5HT7R:::ant::D|||
Ornidazole|inv||||
Biapenem|inv||||
Fenoverine|inv||||
Tirilazad|inv|5HT2C::::6.42:C;5HT2A::::6.24:C;FYN::::5.95:C;ADA2C::::5.94:C;MK14::::5.13:C|||
Parthenolide|ok_inv|PGH2::::6.1:C;NOS2::MOUSE::5.98:C;NFKB2::::5.47:C|||
Tramazoline|inv|ADA2C::RAT::8.38:C;ADA1B::RAT::5.96:C|||
Nimustine|inv|NFKB1::::7.4:C;LMNA::::5.65:C|||
Creatinolfosfate|inv||||
Macimorelin|ok_inv|GHSR:::ago:7.64:DC|CP3A4:::sub::D||
Yttrium_Y_90|ok_inv||||
Pyritinol|inv||||
Riamet|ok_inv||||
Enoxolone|inv|DHI2::::8.92:C;DHI1::MOUSE::8.7:C;DHI1::::8.07:C;LMNA::::7.05:C;DHI1::RAT::7.05:C;KPCL::::6.6:C;SO1B1::::6.54:C;DHI2::RAT::6.44:C;SO1B3::::6.38:C;AK1BA::::5.31:C;PTN11::::5.02:C;CYSP::TRYCR::5.:C|||
Tiropramide|inv||||
Meclocycline|inv|RS7::ECOLI:ant::D|TETX::BACT4:sub::D|OMPF::ECOLI:sub::D;Membrane_protein::ECOLX:sub::D|
Valnoctamide|inv||||
Biguanide|ok_inv||||
Amitriptylinoxide|ok_inv|CP2CJ::::6.4:C;CP1A2::::6.1:C;CP3A4::::5.9:C;RET::::5.:C|||
Norflurane|ok_exp||||
Pentafluoropropane|ok_inv||||
Troxerutin|inv||||
Lusutrombopag|ok_inv|TPOR:::ago::D|CP4AB:::sub::D|MDR1:::inh::D;ABCG2:::sub::D|
Trimegestone|inv||||
Artemisinin|inv||CP2B6:::sub_ind::D||
Von_Willebrand_Factor_Human|ok_inv|FA8:::stbz::D;CO1A1:::bin::D|ATS13:::sub::D||
Fluindione|ok_inv|LOX5::RAT::5.02:C|CP3A4:::sub::D;CP2C9:::sub::D||
Levosalbutamol|ok_inv|HIF1A::::8.49:C;TSHR::::6.9:C;ADRB2:::ago:6.84:DC;NFKB1::::5.2:C|CP2D6:::inh:5.9:DC;CP3A4:::inh::D|SO1B3:::sub::D;SO1B1:::sub::D|
Bezlotoxumab|ok_inv|TOXB::CLODI:abo::D|||
Calcium_glubionate_anhydrous|ok||||
Methallenestril|exp||||
Lenograstim|ok_inv|CSF3R:::ago::D|||
Nedaplatin|ok_inv|Glutathione:::lig::D;DNA:::lig::D|||
Fluciclovine_18F|ok|AAAT:::bin::D;YLAT1:::bin::D;CTR3:::bin::D;NMDA:::inh::D;GRIA1:::inh::D;GRIA2:::inh::D;GRIA3:::inh::D;GRIA4:::inh::D||MDR1:::sub::D;MRP4:::sub::D|
Pancrelipase_lipase|ok|Dietary_fat:::cli::D|||
Coagulation_factor_X_human|ok_inv||||
Protein_S_human|ok|FA5:::ant::D;FA10:::ant::D;PROC:::cof::D|||
Coagulation_factor_VII_human|ok_inv|TF:::act::D;FA10:::act::D;FA9:::act::D|||
Anti_inhibitor_coagulant_complex|ok_inv|FA10:::ago::D;THRB:::ago::D;FIBA:::cli::D;FIBB:::cli::D;F13A:::ago::D;FA5:::ago::D;FA8:::ago::D;FA7:::ago::D|THRB:::sub::D;FA7:::sub::D;FA8:::sub::D;FA9:::sub::D;FA5:::sub::D||
Coagulation_Factor_IX_Human|ok|FA10:::act::D;FA11:::lig::D;FA7:::lig::D;FA8:::cof::D;THRB;LRP1;VKGC|||
Levomenol|ok_exp|||SO1B3:::sub::D;SO1B1:::sub::D|
Parachlorophenol|ok|SCN4A||SO1B3:::sub::D|
Esculin|ok|AL1A1::::6.15:C;PGDH::::5.8:C;CASP7::::5.4:C;CASP1::::5.4:C;CYSP::TRYCR::5.1:C;HCD2::::5.1:C;IMPA1::RAT::5.:C;ANDR:::ago::D|GLSK:::sub::D||
Inosine_pranobex|ok||||
Sodium_lauryl_sulfoacetate|ok_exp||||
Clobetasone|ok|GCR:::ago::D|CP3A4:::sub::D||
Nusinersen|ok_inv|Survival_motor_neuron_protein:::oli::D|EXO::LAMBD:sub::D||
Terpin_hydrate|ok_exp||||
Olmutinib|inv|EGFR:::inh::D|||
Zofenopril|ok|ACE:::inh:9.4:DC|||
Alclofenac|ok_out|PGH2:::ant::D|||
Nandrolone|exp_inv|ANDR::RAT::8.68:C;SHBG::::6.3:C;CBG::::6.14:C|||
Plecanatide|ok_inv|GCYA2:::ago::D|||
Cerliponase_alfa|ok_inv|MPRI:::lig::D|||
Inositol|ok_out|LMNA::::5.:C||SC5A3:::sub::D|
Troleandomycin|ok|NR1I2:::act::D;RL4::ECOLI:inh::D;RL32::DEIRA:inh::D|CP3A4:::inh:5.1:DC;CP3A7:::inh::D;CP2C8:::inh::D;CP343:::ind::D;CP3A5:::inh::D|MDR1:::inh::D|
Gluconic_Acid|ok_inv||||
Technetium_Tc_99m_etifenin|exp||||
Oxabolone_cipionate|exp||||
Calcitonin_porcine|exp||||
Phosphocreatine|nutra|GAMT:::pro::D;SC6A8;KCRM:::lig::D;KCRU:::lig::D;KCRS:::lig::D;KCRB:::lig::D|||
Antihemophilic_factor_human|ok|FA9:::act::D;FA10:::act::D|PROC:::sub::D||
Vitex_agnus_castus_fruit_extract|exp||||
Hedera_helix_leaf_extract|exp||||
Horse_chestnut|exp||||
Valerian|ok_exp_inv||||
Kallidinogenase|exp||||
Pepsin|ok_exp_inv||||
Brinase|exp||||
Lipegfilgrastim|ok_inv|CSF3R:::ago::D|||
Piprozolin|exp||||
Bamifylline|exp||CP1A2:::sub::D||
Dimethyl_carbate|exp||||
Teclozan|exp||||
Bamethan|exp||||
Arginine_glutamate|inv||||
Prednylidene|exp||CP3A4:::sub_ind::D;CP3A5:::ind::D||
Bismuth_subnitrate|ok||||
Sodium_chlorite|exp||||
Guanoxan|ok||||
Phenolsulfonphthalein|exp||||
Butaperazine|ok||||
Sulfadicramide|exp||||
Sulfobromophthalein|exp||||
Oxolamine|ok||||
Fentiazac|exp|PD2R2::::6.26:C|||
Mandelic_acid|ok||||
Medifoxamine|ok||||
Ferrous_aspartate|exp||||
Apronalide|ok||||
Tilbroquinol|ok||||
Fluocortin|exp||||
Piperidione|exp||||
Dibenzepin|ok||||
Acetylleucine|exp||||
Tribenoside|exp||||
Flosequinan|ok||||
Enibomal|exp||||
Gestonorone|exp||||
Calcium_lactate|ok_inv_vet||||
Suxibuzone|exp||||
Alaproclate|exp|SC6A4::RAT::6.15:C|||
Propanidid|exp||||
Perboric_acid|ok||||
Stibophen|exp||||
Clofoctol|exp||||
Tuaminoheptane|exp||||
Neltenexine|exp||||
Cymarin|exp||||
Begelomab|exp_inv||||
Bucladesine|exp||||
Tiazofurine|exp||||
Aminomethylbenzoic_acid|exp||||
Thiram|ok_exp||||
Quinupramine|ok||||
Pramiracetam|ok||||
Phthalylsulfathiazole|ok||||
Magnesium_silicate|ok||||
Methylmethionine_chloride|exp||||
Octopamine|exp||||
Tropatepine|exp||||
Proxibarbal|ok||||
Prifinium|exp||||
Propatyl_nitrate|exp_inv||||
Clothiapine|ok||||
Ferrous_sulfate_anhydrous|ok|Free_radicals:::ago::D|NDUS8;SDHA:::lig::D;XDH:::lig::D;ACON:::cof::D;CP4AB:::cof::D;SUOX:::cof::D;PERM:::lig::D;CATA:::lig::D;NOS2:::lig::D;PGH1:::lig::D;PGH2:::lig::D;TPH1:::lig::D;P4HA1:::lig::D;PHS:::lig::D;CERU:::sub::D|TRFE:::tra::D;FRIL:::sto::D;FRIH:::sto::D;B2ZDZ3:::tra::D;Iron_ABC_transporter_substrate_binding_protein::MANHA:tra::D|
Etofamide|ok||||
Ethyl_chloride|ok_exp_inv||||
Lysozyme|exp_inv||||
Sitafloxacin|exp_inv||CP1A2:::inh::D||
Aceclidine|ok||||
Quassia|exp||||
Penimepicycline|exp||||
Hexobendine|ok||||
Cefatrizine|exp||||
Ritiometan|ok||||
Acetarsol|ok_out||||
Dichlorobenzyl_alcohol|ok|SCN1A:::ant::D|||
Dibekacin|ok||||
Wood_creosote|exp_inv||||
Meladrazine|exp||||
Sultopride|ok||||
Micronomicin|ok||||
Clorindione|exp||CP3A4:::sub::D||
Idanpramine|exp||||
Benziodarone|ok_out||||
Bucetin|ok_out||||
Carbocromen|ok_out||||
Aluminium_acetoacetate|exp||||
Bromelains|inv||||
Benzododecinium|ok||||
Sulfaisodimidine|exp||||
Meticrane|ok||||
Etilamfetamine|exp||||
Bumadizone|ok||||
Miocamycin|ok||CP3A4:::inh::D||
Tromantadine|ok||||
Rimazolium|exp||||
Olaflur|exp||||
Cloridarol|exp||||
Pimethixene|ok||||
Ipecac|ok_out||CP2D6:::sub::D;CP3A4:::sub::D||
Azidamfenicol|exp||||
Atracurium|ok_exp_inv||||
Propamidine|exp_inv|ACRO::PIG::5.46:C;NMDZ1::RAT::5.26:C|||
Idrocilamide|exp||||
Alsactide|exp||||
Sulglicotide|exp||||
Epicillin|exp||||
Hachimycin|exp||||
Febarbamate|exp||||
Triaziquone|exp||||
Tolpropamine|exp||||
Chlorquinaldol|ok||||
Proscillaridin|exp||||
Oxametacin|exp||||
Benproperine|exp||||
Ormeloxifene|exp||||
Trepibutone|exp||||
Delapril|inv||||
Melevodopa|exp||||
Alminoprofen|exp||||
Sobrerol|exp||||
Ibopamine|exp||||
Flunoxaprofen|exp||||
Demecolcine|exp||||
Propenidazole|exp||||
Sulfaperin|exp||||
Methiodal|exp||||
Hydrotalcite|ok_exp_inv||||
Trichloroethylene|ok|TSHR::::8.4:C|||
Tetrazepam|exp||||
Nifurzide|exp||||
Euflavine|exp||||
Picotamide|exp||||
Butanilicaine|exp||||
Guaiazulen|exp||||
Amezinium_metilsulfate|exp||||
Pyrithyldione|exp||||
Dibutylsuccinate|exp||||
Efloxate|exp||||
Mannosulfan|exp||||
Pinazepam|exp||||
Dimethylphthalate|exp||||
Pheneticillin|ok||||
Flurithromycin|exp||CP3A4:::inh::D||
Etoglucid|exp||||
Suloctidil|exp||||
Fenozolone|exp||||
Cinepazet|exp||||
Tioxolone|exp||||
Mercuric_amidochloride|exp||||
Dihydroergocristine|ok_exp|5HT1A:::ant::D;ADRB1:::duo::D;ADA1A:::duo::D;DRD1:::duo::D|CP3A4:::sub::D|ABCBB:::sub::D|
Bufexamac|ok_out|LOX5::RAT::6.89:C;CP1A2::::5.8:C;HIF1A::::5.1:C;FRIL::HORSE::5.05:C;CP2D6::::5.:C;HDA10:::inh::D;HDAC6:::inh::D;PGH2:::inh::D;PGH1:::inh::D|||
Diphenadione|exp||CP3A4:::sub::D||
Tiadenol|exp||||
Talastine|exp||||
Azanidazole|exp||||
Piperidolate|exp||||
Deanol|exp||||
Viminol|exp||||
Phenprobamate|exp||||
Visnadine|exp_inv||||
Mesulfen|exp||||
Styramate|exp||||
Cibenzoline|exp||||
Magnesium_aspartate|exp||||
Tolciclate|exp||||
Trimethyldiphenylpropylamine|exp||||
Pheneturide|exp||||
Oxaceprol|exp||||
Feprazone|exp||||
Calcium_lactate_gluconate|exp||||
Hydrochloric_acid|exp||||
Cloricromen|exp||||
Motretinide|exp||||
Benzilone|exp||||
Bromisoval|exp||||
Difenpiramide|exp||||
Calcium_alginate|ok_exp||||
Acriflavinium_chloride|exp||||
Vincamine|exp||||
Edrecolomab|exp_inv||||
Succinimide|exp||||
Vinbarbital|exp||||
Norfenefrine|exp||||
Chiniofon|exp||||
Difemerine|exp||||
Sodium_feredetate|ok||||
Chlorproethazine|exp||||
Diiodohydroxypropane|exp||||
Melitracen|exp_inv||||
Dihydroergocryptine|exp||CP3A4:::sub::D||
Epimestrol|exp||||
Hematin|exp||||
Phenylmercuric_nitrate|exp||||
Iopydol|exp||||
Levoverbenone|exp||||
Mercurochrome|exp||||
Emetine|exp||||
Adrenalone|exp||||
Eprozinol|exp||||
Neocitrullamon|exp||||THBG:::sub::D
Prenoxdiazine|exp||||
Oxyfedrine|exp||||
Terguride|exp||CP3A4:::sub::D||
Linsidomine|exp||||
Metildigoxin|exp||||
Acetylglycinamide_chloral_hydrate|exp||||
Oxypertine|exp||||
Edetate_sodium|exp||||
Mefruside|exp||||
Carbutamide|exp||CP2C9:::sub::D||
Nifenazone|exp||||
Methylpropylpropanediol_dinitrate|exp||||
Rokitamycin|exp||CP3A4:::inh::D||
Guanoxabenz|exp||||
Lofepramine|exp||||
Pirisudanol|exp||||
Phenglutarimide|exp||||
Fenyramidol|exp||||
Pentetrazol|exp||||
Sulbutiamine|exp||||
Morinamide|exp||||
Moxestrol|exp||||
Troxipide|exp||||
Thiazinam|exp||||
Edoxudine|ok_out|LMNA::::6.35:C;DNA_polymerase::HHV1:inh::D|||ALBU:::bin::D
Nicofuranose|exp||||
Ferric_hydroxide|exp||||
Clofenotane|exp||||
Flutrimazole|exp||||
Gold_Au_198|exp||||
Iobenzamic_acid|exp||||
Tolonidine|exp||||
Mebutizide|exp||||
Proglumide|exp||||
Lonazolac|exp||||
Simfibrate|exp||||
Fenticonazole|exp||||
Endralazine|exp||||
Droxypropine|exp||||
Medazepam|exp||||
Prolintane|exp||||
Fenpiprane|exp||||
Niceritrol|exp||||
Citiolone|exp||||
Esatenolol|exp||CP2D6:::sub::D||
Ioxitalamic_acid|ok_exp||||
Nepinalone|exp||||
Guar_gum|exp||||
Prethcamide|exp||||
Mazaticol|exp||||
Proxyphylline|exp||CP1A2:::sub::D||
Tioclomarol|exp||||
Cadralazine|exp||||
Xenon|exp||||
Nicomorphine|exp||||
Phenibut|exp||||
Midecamycin|exp||CP3A4:::inh::D||
Oxaflozane|exp||||
Thebacon|exp||||
Pecilocin|exp||||
Ronifibrate|exp||||
Cefcapene|exp||||
Bephenium|exp||||
Oxetorone|exp||||
Ornipressin|exp||||
Ciclobendazole|exp||||
Deptropine|exp||||
Lanatoside_C|exp||||
Etybenzatropine|exp||||
Phanquinone|exp||||
Cefodizime|exp||||
Nalfurafine|exp_inv|OPRK::::10.6:C;OPRK::CAVPO::9.77:C;OPRD::RAT::9.43:C;OPRM::CAVPO::9.41:C;OPRM::MOUSE::9.37:C;OPRM::::9.14:C;OPRD::MOUSE::7.29:C;OPRD::::7.13:C|||
Cyclofenil|exp||||
Antimony_pentasulfide|exp||||
Tipepidine|exp||||
Furazidin|exp||||
Diisopromine|exp||||
Sodium_apolate|exp||||
Meptazinol|exp||||
Histapyrrodine|exp||||
Lentinan|exp_inv||||
Tenidap|exp||||
Dimefline|exp||||
Etamsylate|exp||||
Quinbolone|exp||||
Sulfametomidine|exp||||
Magnesium_peroxide|exp||||
Iodine_131I_norcholesterol|exp||||
Bencyclane|exp||CP3A4:::sub::D||
Bamipine|exp||||
Hidrosmin|exp||||
Fluperolone|exp||||
Policresulen|exp_inv||||
Cyclobutyrol|exp||||
Dimetofrine|exp||||
Paraoxon|exp||||
Iprindole|exp||||
Valethamate|exp||||
Cefsulodin|exp||||
Otilonium|exp_inv||CP3A4:::sub::D||
Bendazac|ok_out|Free_radicals:::inh::D;PGH1;PGH2|||
Budipine|exp||||
Tyrothricin|ok|ACES:::inh::D;BGAL::ECOLI:inh::D;Phospholipid_membrane::ECOLI:disrupt::D|||
Cefetamet|exp||||
Emepronium|exp||||
Carfecillin|exp||||
Poldine|exp||||
Cloranolol|exp||CP2D6:::sub::D||
Aloxiprin|exp||||
Buflomedil|exp||||
Clebopride|exp||||
Clefamide|exp||||
Tribromometacresol|exp||||
Pranoprofen|exp_inv|PGH1::RAT::6.41:C;PGH1::SHEEP::5.51:C|||
Levomethadone|exp||||
Clodantoin|exp||||
Angiotensinamide|exp||||
Alginic_acid|ok_inv||||
Cerium_oxalate|exp||||
Metergoline|ok|5HT2A::::9.95:C;5HT2B::::9.55:C;5HT2B::RAT::9.52:C;5HT2C::::9.46:C;5HT1A::::8.64:C;DRD3::::8.58:C;5HT1A::RAT::8.45:C;5HT7R::::8.2:C;5HT7R::RAT::8.2:C;ADA2B::::8.12:C;5HT1B::RAT::7.96:C;5HT6R::::7.89:C;DRD2::::7.68:C;ADA2A::::7.66:C;ADA2C::::7.57:C;DRD1::::7.43:C;ADA1A::RAT::7.42:C;SC6A3::::7.3:C;ADA1D::::7.17:C;ADA1B::RAT::6.84:C;CP2D6::::6.7:C;5HT4R::CAVPO::6.56:C;SC6A4::::6.5:C;SC6A2::::6.44:C;HRH1::::6.32:C;HRH2::::6.02:C;TAU::::6.:C;ACES::::5.87:C;NK2R::::5.87:C;MEN1::::5.6:C;LMNA::::5.15:C;UBP2::::5.:C;TPO::::5.:C;SCN2A:::inh::D|||
Alipogene_tiparvovec|ok_inv||||
Mebicar|exp||||
Veralipride|exp||||
Propyphenazone|exp||||
Althea_root|exp||||
Pentaerithrityl|exp||||
Proglumetacin|exp||||
Chlormadinone|exp||CP3A4:::sub::D||
Dobesilic_acid|exp_inv||||
Mepindolol|exp||CP2D6:::sub::D||
Nicofetamide|exp||||
Cyclopenthiazide|ok||||
Methylestrenolone|exp||||
Gedocarnil|exp||||
Nebacumab|exp||||
Broxyquinoline|exp||||
Gitoformate|exp||||
Guacetisal|exp||||
Iodoxamic_acid|exp||||
Isepamicin|exp||||
Iprazochrome|exp||||
Bevonium|exp||||
Mitobronitol|exp||||
Ethenzamide|exp||||
Isobromindione|exp||||
Nizofenone|exp||||
Sulfatolamide|exp||||
Dibrompropamidine|exp||||
4_dimethylaminophenol|exp||||
Bifemelane|exp||||
Cinchophen|exp||||
Trifluperidol|exp||||
Carumonam|exp||||
Moperone|exp||||
Prajmaline|exp||||
Sulfamazone|exp||||
Thiopropazate|exp||||
Morclofone|exp||||
Rimiterol|exp||||
Dextranomer|exp||||
Clobenzorex|exp||||
Norgestrienone|exp||||
Zipeprol|exp||||
Benzoxonium|exp||||
Sequifenadine|exp||||
Desaspidin|exp||||
Diodone|exp||||
Ferrous_chloride|exp||||
Oxidized_cellulose|exp||||
Pentamycin|exp||||
Emylcamate|exp||||
Acefylline|exp||CP1A2:::sub::D||
Heptaminol|exp||||
Bietaserpine|exp||||
Aluminium_nicotinate|exp||||
Allobarbital|exp||||
Metabutethamine|exp||||
Mepixanox|exp||||
Succinylsulfathiazole|exp||||
Rociverine|exp|ACM1:::ant::D;ACM2:::ant::D;ACM3:::ant::D;ACM4:::ant::D;ACM5:::ant::D|||
Ferric_59Fe_citrate|exp||||
Mephenesin|ok||||
Gallamine|exp||||
Aminoethyl_nitrate|exp||||
Metandienone|exp||||
Mesterolone|exp|SHBG::::9.6:C|||
Naftidrofuryl|exp||||
Calcium_pangamate|exp||||
Metopimazine|exp||||
Etamiphylline|exp||CP1A2:::sub::D||
Zolimidine|exp||||
Almasilate|ok_exp||||
Oxycinchophen|exp||||
Moroxydine|exp||||
Diethyl_ether|exp||||
Difetarsone|exp||||
Deltamethrin|exp||||
Oxiracetam|exp||||
Promegestone|exp||CP3A4:::sub::D||
Pyrrolnitrin|exp||||
Guanazodine|exp||||
Phenoperidine|exp||||
Phenazocine|exp||||
Picloxydine|exp||||
Tiocarlide|exp||||
Umifenovir|exp_inv|LYAG::::5.05:C|||
Flumedroxone|exp||||
Chlormidazole|exp||||
Carbaspirin_calcium|exp_inv||||
Ticlatone|exp||||
Metizoline|exp||||
Mifamurtide|ok_exp|TLR4:::lig::D;NOD2:::lig::D|||
Melagatran|exp||||
Clorexolone|exp||||
Ipriflavone|exp||||
Bornaprine|exp||||
Potassium_gluconate|ok||ATNG:::sub_ind::D|AT1A1:::sub::D;S12A1:::sub::D;ATP4A:::sub::D|
Tetragalacturonic_acid_hydroxymethylester|exp||||
Selenium_75Se_norcholesterol|exp||||
Fabomotizole|exp||||
Methoxyphenamine|ok||||
Carbuterol|exp||||
Aluminium_glycinate|exp||||
Oxolinic_acid|exp||CP1A2:::inh::D||
Ethyl_hydroxybenzoate|ok_exp||||
Mofebutazone|exp||||
Bibenzonium|exp||||
Methoserpidine|exp||||
Protiofate|exp||||
Mepartricin|exp||CP3A4:::inh::D||
Pentifylline|exp||CP1A2:::sub::D||
Tiracizine|exp||||
Etanautine|exp||||
Tenitramine|exp||||
Cefbuperazone|exp||||
Ferrous_tartrate|exp||||
Acetoxolone|exp||||
Metisazone|exp||||
Pridinol|exp||||
Loprazolam|exp||||
Methylthiouracil|exp||||
Ethacizine|exp||||
Saruplase|exp||||
Semustine|exp_inv||||
Alcuronium|exp||||
Proquazone|exp||||
Aloglutamol|exp||||
Lorajmine|exp||||
Bunaftine|exp||||
Lorcainide|exp||||
Montmorillonite|exp_inv||||
Nikethamide|exp||||
Eberconazole|exp||||
Benorilate|ok||||
Hemoglobin_raffimer|exp_inv||||
Tenonitrozole|exp||||
Propicillin|exp||||
Niridazole|exp||||
Hexapropymate|exp||||
Clofenamide|exp||||
Formocortal|exp||||
Fluanisone|exp||||
Tiemonium_iodide|exp||||
Cefozopran|exp||||
Ipidacrine|exp||||
Morpholine|exp||||
Oxantel|exp||||
Sulbentine|exp||||
Dimethylaminopropionylphenothiazine|exp||||
Bekanamycin|exp||||
Cridanimod|exp||||
Metahexamide|exp||CP2C9:::sub::D||
Mosapramine|exp||||
Carboquone|exp||||
Dihexyverine|exp||||
Dexchlorpheniramine|exp_inv|HRH1::::9.14:C;SC6A4::::7.89:C;ACM4::::6.56:C;ACM1::::6.48:C;ACM3::::6.26:C;SGMR1::::6.16:C;SC6A3::::6.13:C;ACM5::::6.13:C;5HT2A::::5.98:C;5HT2C::::5.91:C;ADA2B::::5.68:C;ACM2::::5.6:C;SC6A2::::5.31:C;ADA2A::::5.12:C;HRH2::::5.08:C;ADA1B::RAT::5.06:C|CP2D6:::inh::D||
Naftazone|ok||||
Butalamine|exp||||
Cefpirome|ok||||
Quinisocaine|exp||||
Omoconazole|exp||||
Quingestanol|exp||CP3A4:::sub::D||
Clometocillin|exp||||
Niaprazine|exp||||
Drisapersen|exp_inv||||
Tacalcitol|exp_inv|VDR::::8.15:C|||
Vinyl_ether|exp||||
Acetyldigoxin|exp||||
Tretoquinol|exp||||
Sulbenicillin|exp||||
Distigmine|exp||||
Penthienate|exp||||
Bromochlorosalicylanilide|exp||||
Ambazone|exp||||
Ferrous_carbonate|exp||||
Sulfathiourea|exp||||
Protamine|exp_inv||||
Ioglicic_acid|exp||||
Tibezonium_iodide|exp||||
Gepefrine|exp||||
Pristinamycin|exp_inv||||
Decamethoxine|exp||||
Eosin|exp||||
Sodium_tartrate|ok||||
Fenquizone|exp||||
Ciclonicate|exp||||
Metenolone|exp||||
Tritoqualine|ok||||
Dixanthogen|exp||||
Quifenadine|exp||||
Xibornol|exp||||
Dilazep|exp||||
Dibutylphthalate|exp||||
Phenothrin|exp||||
Hydroquinine|exp||||
Trolnitrate|exp||||
Diphemanil|ok_vet_out|ACM3:::ant::D|||
Cypermethrin|exp||||
Pirprofen|exp||||
Meldonium|exp||||
Nifuratel|exp||||
Terodiline|exp||CP3A4:::sub::D||
Sulfaguanidine|exp||||
Azapetine|exp||||
Halometasone|exp||CP3A4:::ind::D;CP3A5:::ind::D||
Camostat|exp||||
Nifurtoinol|exp||||
Butamirate|exp||||
Meglumine_antimoniate|exp_inv||||
Methylpentynol|exp||||
Biphenylol|exp||||
Fenoxazoline|exp||||
Cyclobarbital|exp||||
Camylofin|exp||||
Penamecillin|exp||||
Bemegride|exp||||
Ioglycamic_acid|exp||||
Elcatonin|exp||||
Sodium_aurotiosulfate|ok_exp||||
Piromidic_acid|exp||||
Fazadinium_bromide|exp||||
Bioallethrin|ok_exp|SCN1A:::mod::D;Sodium_channel_protein::9NEOP:mod::D;CCG1:::ago::D;CAC1G:::inh::D;CAC1A:::inh::D;CAC1C:::inh::D|CP2C8:::sub::D;CP2C9:::sub::D;CP2CJ:::sub::D;CP3A4:::sub::D;CP2A1::RAT:sub::D;CP1A1::RAT:sub::D;CP2C6::RAT:sub::D;CP2CB::RAT:sub::D;CP3A1::RAT:sub::D;CP3A2::RAT:sub::D||
Trolamine|ok||||
Tidiacic_arginine|exp||||
Magnesium_gluconate|ok_inv||HXK::SCHMA:sub::D;KCRB:::sub_ind::D;ABL1:::sub_ind::D;ATPD:::sub::D;ADCY1:::sub::D;GCYA2:::sub::D;F261:::ind::D;Phosphoribosylpyrophosphate_synthetase::PLAF7:ind::D;AT1A1:::ind::D||
Obidoxime|exp||||
Glycyrrhizic_acid|ok_exp|DHI1:::ant::D;TNFA:::ant::D;CASP3:::ant::D;NFKB2:::inh::D;LIPL:::ind::D||ABCBB:::sub::D|AK1C4:::sub::D;AK1C3:::sub::D;AK1C2:::sub::D;ALBU:::sub::D
Tetramethrin|exp||||
Cetiedil|exp||||
Mephenoxalone|exp||||
Iocarmic_acid|exp||||
Peruvoside|exp||||
Epanolol|exp||CP2D6:::sub::D||
Meclofenoxate|exp||||
Fenpiverinium|exp||||
Niperotidine|exp_inv||||
Tilactase|ok_exp|Lactose:::cli::D|||
Dexrabeprazole|exp||CP2CJ:::sub::D||
Aurotioprol|exp||||
Monoxerutin|exp||||
Mercuric_chloride|exp||||
Lidoflazine|ok_exp||CP3A4:::sub::D||
Vorozole|exp||||
Domiodol|exp||||
Emetonium_iodide|exp||||
Vinylbital|exp||||
Ferric_sodium_citrate|exp||||
Rufloxacin|exp|MK01::::5.2:C|CP1A2:::inh::D||
Sulfamethoxypyridazine|exp||||
Myristalkonium|exp||||
Tertatolol|exp||CP2D6:::sub::D||
Ibacitabine|exp||||
Prenalterol|exp||||
Cefazedone|exp||||
Guanoclor|exp||||
Aluminium_clofibrate|exp||||
Xamoterol|ok_exp|ADRB1:::pag:7.96:DC;ADRB2::::6.18:C|||
Imipramine_oxide|exp||||
Acemetacin|ok_inv|HIF1A::::7.:C;PGH2:::ant::D;PGH1:::ant::D|UD2B7:::sub::D|MRP1:::sub::D|
Dixyrazine|exp||||
Dropropizine|exp||||
Magnesium_orotate|exp||||
Tilidine|exp||||
Chlorbenzoxamine|exp||||
Aluminium_acetotartrate|exp||||
Fipexide|exp||||
Penfluridol|exp||CP3A4:::sub::D||
Clopamide|exp|LMNA::::6.5:C|||
Vinburnine|exp||||
Dimethoxanate|exp||||
Brodimoprim|exp||||
Dibunate|exp||||
Iodocholesterol_131I|exp||||
Demoxytocin|exp||||
Ethadione|exp||||
Calcium_levulinate|ok_exp|CALM1:::ago::D;CASQ1:::ago::D;CALB2:::ago::D|||
Muzolimine|ok_out||||
Epomediol|exp||||
Xipamide|exp||||
Benzylthiouracil|exp||||
Reposal|exp||||
Linopirdine|exp||||
Tisopurine|exp||||
Mebhydrolin|exp||||
Paclitaxel_poliglumex|exp_inv||||
Dimemorfan|exp||||
Oblimersen|exp_inv||||
Bufylline|exp||CP1A2:::sub::D||
Iodoform|ok_exp_vet||||
Talampicillin|exp||||
Xenysalate|exp||||
Aspoxicillin|exp||||
Carbromal|exp||||
Bibrocathol|exp||||
Proxazole|exp||||
Oxomemazine|exp||||
Ceftezole|exp||||
Meprotixol|exp||||
Pipemidic_acid|exp||CP1A2:::inh::D||
Enprostil|exp||||
Fedrilate|exp||||
Etohexadiol|exp||||
Indanazoline|exp||||
Cyfluthrin|exp||||
Calcium_silicate|exp||||
Copper_usnate|exp||||
Potassium_permanganate|exp_inv||||
Ranimustine|exp||||
Methylatropine|exp||||
Phenylmercuric_borate|exp||||
Caroverine|exp||CP3A4:::sub::D||
Metampicillin|exp||||
Doxefazepam|exp||||
Noxytiolin|ok||||
Dipyrocetyl|exp||||
Hydroxyethylpromethazine|exp||||
Clopenthixol|exp||||
Etofylline_nicotinate|exp||||
Cloprednol|exp||CP3A4:::ind::D;CP3A5:::ind::D||
Pipenzolate|exp||||
Etafenone|exp||||
Pyrrobutamine|exp||||
Rhenium_Re_186_sulfide|exp||||
Fluorodopa_18F|ok_exp||||
Clofibride|exp||||
Timepidium|exp||||
Artemotil|ok||||
Mefenorex|exp||||
Anethole_trithione|ok_exp||||
Gamolenic_acid|ok_inv|PPARA::::6.57:C;CASP6::::6.3:C;PPARD::::6.12:C;PPARG::::5.66:C;FFAR1::::5.34:C;AMPC::ECOLI::5.3:C|||
Nifuroxazide|exp||||
Fluclorolone|exp||||
Demegestone|exp|PRGR:::ago::D|CP3A4:::sub::D||
Dimazole|ok_out|LMNA::::5.85:C|||
Imidazole_salicylate|exp||||
Iopentol|exp||||
Magnesium_phosphate|exp||||
Fosfructose|exp|KPYM::::7.64:C;ALF::TRYBB::5.:C|||
Hemoglobin_crosfumaril|exp||||
Dehydroemetine|inv||||
Etynodiol|exp||CP3A4:::sub::D||
Fluticasone|ok_exp|GCR:::ago::D;PRGR:::ago::D;PA24A:::inh::D;MCR:::ant::D|CP3A4:::duo::D;CP3A5:::duo::D;CP3A7:::sub::D;CP2C8:::inh::D|MDR1:::sub::D;SO1B1:::inh::D|CBG;MDR1:::sub::D;SO1B1:::inh::D
Lormetazepam|ok|GBRA2:::aga::D;GBRG2:::aga::D;GBRA3:::aga::D;GBRA5:::aga::D;GBRA1:::aga::D|||
Fenofibric_acid|ok|FABPL::RAT::7.03:C;FABPI::::6.:C;PPARA:::ago:5.58:DC;NR1I2:::pag::D;PPARD;PPARG;MMP25|||
Enasidenib|ok_inv|IDHP:::inh::D|CP1A2:::inh::D;CP2B6:::duo::D;CP2C8:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D;CP2D6:::inh::D;CP3A4:::duo::D;UD11:::inh::D;UD13:::sub::D;UD14:::sub::D;UD19:::sub::D;UD2B7:::sub::D;UDB15:::sub::D|MDR1:::inh::D;ABCG2:::inh::D;S22A6:::inh::D;SO1B1:::inh::D;S22A2:::inh::D;SO1B3:::inh::D;S22A8:::inh::D|
Pibrentasvir|ok_inv|Nonstructural_protein_5A::9HEPC:inh::D|CP3A4:::inh::D;UD11:::inh::D|MDR1:::inh::D;ABCG2:::inh::D;SO1B1:::inh::D;SO1B3:::inh::D|
Glecaprevir|ok_inv|NS3_protease::9HEPC:inh::D|CP3A4:::inh::D;UD11:::inh::D;CP3A4:::inh::D|MDR1:::inh::D;ABCG2:::inh::D;SO1B1:::inh::D;SO1B3:::inh::D|
Tisagenlecleucel|ok_inv|CD19:::abo::D|||
Methyl_nicotinate|ok|AL1A1::::7.6:C|||
Coral_snake_micrurus_fulvius_immune_globulin_antivenin_equine|ok_exp||||
Albutrepenonacog_alfa|ok|FA10:::act::D|FA8:::sub::D||
Ferric_subsulfate|ok_exp||||
Human_cytomegalovirus_immune_globulin|ok||||
Meningococcal_polysaccharide_vaccine_group_W_135|ok_exp_inv||||
Meningococcal_polysaccharide_vaccine_group_Y|ok_exp_inv||||
Meningococcal_polysaccharide_vaccine_group_A|ok_exp_inv||||
Meningococcal_polysaccharide_vaccine_group_C|ok_exp_inv||||
Crotalus_scutulatus_antivenin|ok_exp||||
Crotalus_atrox_antivenin|ok_exp||PA2GX:::inh::D||
Crotalus_adamanteus_antivenin|ok_exp|PA2GX:::ant::D|ENPP1:::lig::D;PA2GX:::inh::D||
Agkistrodon_piscivorus_antivenin|ok_exp|PA2GX:::ant::D|||
Rhus_Glabra_Pollen|ok_exp||||
Talimogene_laherparepvec|ok_exp_inv|Heparan_sulfate;DPOL::HHV11:act::D;DPOL::VZVD:act::D|||
Equine_Botulinum_Neurotoxin_E_Immune_FAB2|ok_exp_inv|BXE::CLOBO:abo::D|||
Equine_Botulinum_Neurotoxin_C_Immune_FAB2|ok_exp_inv|BXC::CBCP:abo::D|||
Equine_Botulinum_Neurotoxin_G_Immune_FAB2|ok_exp_inv|BXG::CLOBO:abo::D|||
Equine_Botulinum_Neurotoxin_A_Immune_FAB2|ok_exp_inv|BXA1::CLOBO:abo::D|||
Equine_Botulinum_Neurotoxin_F_Immune_FAB2|ok_exp_inv|BXF::CLOBO:abo::D|||
Equine_Botulinum_Neurotoxin_D_Immune_FAB2|ok_exp_inv|BXD::CBDP:abo::D|||
Equine_Botulinum_Neurotoxin_B_Immune_FAB2|ok_exp_inv|BXB::CLOBO:abo::D|||
Cat_dander_extract|ok||||
Scorpion_centruroides_immune_Fab2_antivenin_equine|ok||||
Aloe_Vera_Leaf|ok_exp|Free_radicals:::chel::D|||
Fusarium_graminearum|ok_exp||||
Amylmetacresol|ok|SCN2A:::ant::D|||
Bismuth_subgallate|ok||||ALBU:::car::D
Valproate_bismuth|ok||||
Phloxine_B|ok||||
Belladonna|ok_exp||||
Axicabtagene_ciloleucel|ok|CD19:::abo::D|||
Candesartan|exp|AGTR1::RABIT::9.19:C;AGTR1:::ant:9.16:DC;AGTRA::RAT::8.5:C;AGTR1::BOVIN::6.96:C;AA3R::::6.16:C;ADA2B::::5.76:C;SC6A2::::5.52:C;THAS::::5.51:C;ADRB3::::5.49:C;EGFR::::5.48:C;ERBB2::::5.23:C;CP3A4::::5.05:C|CP2C9:::inh:5.52:DC;PGH1:::sub::D;UD13:::sub::D;CP2C8:::inh::D|SO1B1:::inh::D;MDR1:::inh::D|
Emicizumab|ok_inv|FA9:::cof::D;FA10:::act::D|||
Varicella_Zoster_Vaccine_Recombinant|ok_inv||||
Dotatate_gallium_Ga_68|ok_inv|SSR2:::bin::D|||
Cenegermin|ok_inv|NTRK1:::sti::D|||
Semaglutide|ok_inv|GLP1R:::ago::D|DPP4:::sub::D;NEP:::sub::D;LIPL:::inh::D;AMY1:::inh::D||ALBU:::sub::D
Netarsudil|ok|ROCK1:::inh::D;ROCK2:::inh::D;SC6A2:::inh::D|||
Voretigene_neparvovec|ok|RPE65:::gene_replace::D|||
Nonacog_beta_pegol|ok_inv|FA7:::cof::D;FA8:::cof::D;FA10:::ago::D|||
Piperaquine|exp_inv||CP2E1:::ind::D;CP2B6:::inh::D;CP2C9:::sub::D;CP2CJ:::inh::D;CP3A4:::inh::D||
Testosterone_cypionate|ok|ANDR:::ago::D;ESR1;MCR|CP3A4:::duo::D;AOFA:::ind::D;CP11A:::inh::D;CP3A5:::sub::D;CP3A7:::sub::D;CP1A1:::sub::D;CP2AD:::sub::D;CP2B6:::sub_ind::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D;CP343:::sub::D;S5A1:::sub::D;CP19A:::sub::D|SO1A2:::duo::D;S22A8:::ind::D;S22A7:::ind::D;MDR1:::inh::D;NTCP:::inh::D;S22A3:::sub::D;S22A4:::sub::D;ABCG2:::sub::D|ALBU;SHBG
Testosterone_enanthate|ok|ANDR:::ago::D;ESR1;MCR|CP3A4:::duo::D;AOFA:::ind::D;CP11A:::inh::D;CP3A5:::sub::D;CP3A7:::sub::D;CP1A1:::sub::D;CP2AD:::sub::D;CP2B6:::sub_ind::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D;CP343:::sub::D;S5A1:::sub::D;CP19A:::sub::D|SO1A2:::duo::D;S22A8:::ind::D;S22A7:::ind::D;MDR1:::inh::D;NTCP:::inh::D;S22A3:::sub::D;S22A4:::sub::D;ABCG2:::sub::D|ALBU;SHBG
Testosterone_undecanoate|ok_inv|ANDR:::ago::D;ESR1;MCR|CP3A4:::duo::D;AOFA:::ind::D;CP11A:::inh::D;CP3A5:::sub::D;CP3A7:::sub::D;CP1A1:::sub::D;CP1B1:::sub::D;CP2AD:::sub::D;CP2B6:::sub_ind::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D;CP343:::sub::D;S5A1:::sub::D;CP19A:::sub::D|SO1A2:::duo::D;S22A8:::ind::D;S22A7:::ind::D;MDR1:::inh::D;NTCP:::inh::D;S22A4:::sub::D;ABCG2:::sub::D;S22A2;S47A1;SO1B3|ALBU;SHBG
Testosterone_enantate_benzilic_acid_hydrazone|ok_exp||||
Ferric_cation|ok|FHUD::ECOLI:bin::D;TFR1:::ago::D|||TRFE:::bin::D;ITB3:::bin::D;CALR:::bin::D
Estradiol_acetate|ok_inv_vet|ERR3:::lig::D;DHB2;BECN1;ATP6;GPER1;NCOA2;ACHA4;ESR2:::ago::D;NR1I2;ESR1:::ago::D|CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub_ind::D;UD11:::sub::D;CP1A2:::inh::D|SO4A1;SO1C1;SO1B3;S22A8;MDR1:::sub::D;SO1B1:::inh::D;ABCG2:::inh::D;S22AB:::inh::D;MRP7:::inh::D;SO1A2:::inh::D;SO2B1:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|FABPI;ALBU;SHBG
Estradiol_benzoate|ok_inv_vet|ANDR::RAT::8.16:C;ESR1:::ago:7.74:DC;STRP::STRP1::5.72:C;SC6A4::::5.71:C;GCR::::5.64:C;LMNA::::5.5:C;ADA2C::::5.45:C;5HT2B::::5.13:C;ERR3:::lig::D;DHB2;BECN1;ATP6;GPER1;NCOA2;ACHA4;ESR2:::ago::D;NR1I2|CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub_ind::D;UD11:::sub::D;CP1A2:::inh::D|SO4A1;SO1C1;SO1B3;S22A8;MDR1:::sub::D;SO1B1:::inh::D;ABCG2:::inh::D;S22AB:::inh::D;MRP7:::inh::D;SO1A2:::inh::D;SO2B1:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|SHBG::::5.94:DC;FABPI;ALBU
Estradiol_cypionate|ok_inv_vet|ERR3:::lig::D;DHB2;BECN1;ATP6;GPER1;NCOA2;ACHA4;ESR2:::ago::D;NR1I2;ESR1:::ago::D|CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub_ind::D;UD11:::sub::D;CP1A2:::inh::D|SO4A1;SO1C1;SO1B3;S22A8;MDR1:::sub::D;SO1B1:::inh::D;ABCG2:::inh::D;S22AB:::inh::D;MRP7:::inh::D;SO1A2:::inh::D;SO2B1:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|FABPI;ALBU;SHBG
Estradiol_dienanthate|ok_inv_vet|ESR1:::ago::D;NR1I2;ESR2:::ago::D;ACHA4;NCOA2;GPER1;ATP6;BECN1;DHB2;ERR3:::lig::D|CP1A2:::inh::D;UD11:::sub::D;CP3A4:::sub_ind::D;CP3A5:::sub::D;CP3A7:::sub::D;CP1A1:::sub::D;CP1B1:::sub::D;CP2CJ:::sub::D;CP2C8:::sub::D;CP2C9:::sub::D|S22A2:::inh::D;S22A1:::inh::D;S22A3:::inh::D;SO2B1:::inh::D;SO1A2:::inh::D;MRP7:::inh::D;S22AB:::inh::D;ABCG2:::inh::D;SO1B1:::inh::D;MDR1:::sub::D;S22A8;SO1B3;SO1C1;SO4A1|SHBG;ALBU;FABPI
Estradiol_valerate|ok_inv_vet|TAU::::5.8:C;STRP::STRP1::5.42:C;LMNA::::5.25:C;ERR3:::lig::D;DHB2;BECN1;ATP6;GPER1;NCOA2;ACHA4;ESR2:::ago::D;NR1I2;ESR1:::ago::D|CP2C9:::sub::D;CP2C8:::sub::D;CP2CJ:::sub::D;CP1B1:::sub::D;CP1A1:::sub::D;CP3A7:::sub::D;CP3A5:::sub::D;CP3A4:::sub_ind::D;UD11:::sub::D;CP1A2:::inh::D|SO4A1;SO1C1;SO1B3;S22A8;MDR1:::sub::D;SO1B1:::inh::D;ABCG2:::inh::D;S22AB:::inh::D;MRP7:::inh::D;SO1A2:::inh::D;SO2B1:::inh::D;S22A3:::inh::D;S22A1:::inh::D;S22A2:::inh::D|FABPI;ALBU;SHBG
Medium_chain_triglycerides|ok||||
Bronopol|ok|FFP::BACIU::5.05:C;Thiol_groups:::oxi::D|||
Fish_oil|ok_nutra|DGAT2:::ago::D;PGH2:::inh::D;FFAR4:::ago::D;CAC1C:::inh::D;SCN1A:::inh::D;Free_radicals;NFKB2:::reg::D;SRBP1:::reg::D;PPARA:::reg::D;PPARG;PPARD:::reg::D|CP3A4:::sub::D||
Calcium_saccharate|ok_exp||||
Peanut_oil|ok||||
Sarracenia_Purpurea|ok_exp||||
Isopropyl_myristate|ok_exp|LMNA::::6.25:C|||
Patent_Blue|ok|ALBU:::bin::D|||
Plasma_protein_fraction_human|ok||||
Dioctyldimonium|ok_exp||||
Vanadium|ok_exp||||
Racemethionine|ok_exp||||
Remestemcel_L|ok_inv||||
Passiflora_incarnata_flower|ok_exp||||
Black_cohosh|exp||CP3A4:::inh::D;CP3A2::RAT:duo::D;CP1A2:::inh::D;CP2C9:::inh::D;CP2D6:::inh::D||
Sulesomab|ok||||
Potassium_carbonate|ok||||
Besilesomab|ok|Carcinoembryonic_antigen|||
Copper_Cu_64|ok||||
Lutetium_Lu_177|ok||||
Lutetium_Lu_177_dotatate|ok_inv|SSR2:::ago::D;SSR1:::ago::D;SSR3:::ago::D;SSR4:::ago::D;SSR5:::ago::D|||
Strontium_chloride|ok||||
Epitizide|exp||||
Ferric_pyrophosphate_citrate|ok_inv|FRIL:::bin::D;FRIH:::bin::D;HBA:::bin::D;HBB:::bin::D|||
Magnesium_acetate|ok|AT1A1|||
Baloxavir_marboxil|ok_inv|PA::I34A1:inh::D|UD13:::sub::D;CP3A4:::sub::D|ABCB5:::sub::D|
Lonoctocog_alfa|ok_inv|FA10:::act::D;PAHX:::ant::D;FA9:::cof::D;ASGR2:::bin::D;BIP:::chap::D;CALR:::chap::D;CALX:::chap::D;LMAN1:::chap::D;LRP1:::mod::D;MCFD2:::mod::D;VWF:::bin::D|THRB:::act::D;PROC:::inh::D||
Moroctocog_alfa|ok|FA10:::act::D;PAHX:::ant::D;FA9:::cof::D;ASGR2:::bin::D;BIP:::chap::D;CALR:::chap::D;CALX:::chap::D;LMAN1:::chap::D;LRP1:::mod::D;MCFD2:::mod::D;VWF:::bin::D|THRB:::act::D;PROC:::inh::D||
alpha_Tocopherol_succinate|ok_nutra_vet|Lung_epithelial_cells;PP2AA;PP2AB;DGKA;KPCA;LOX5;KPCB;NR1I2;S14L2;S14L3;S14L4|SODC:::ind::D;HMOX1:::ind::D;NQO1:::ind::D;GSH1:::ind::D;GSTM3:::ind::D;GSTO1:::inh::D;GSTP1:::inh::D;GSTA2:::ind::D||TTPA
D_alpha_Tocopherol_acetate|ok_nutra_vet|PP2AA;PP2AB;DGKA;KPCA;LOX5;KPCB;NR1I2;S14L2;S14L3;S14L4|SODC:::ind::D;HMOX1:::ind::D;NQO1:::ind::D;GSH1:::ind::D;GSTM3:::ind::D;GSTO1:::inh::D;GSTP1:::inh::D;GSTA2:::ind::D||TTPA
alpha_Tocopherol_acetate|ok|Free_radicals:::bin::D|CP4F2:::sub::D;CP3A4:::sub::D|TTPA:::sub::D;S14L4:::sub::D;S14L2:::sub::D;S14L3:::sub::D;APOBR:::sub::D;SCRB1:::sub::D;MDR1:::sub::D|VLDLR:::bin::D;LDLR:::bin::D
Tildrakizumab|ok_inv|IL12B:::ant::D|CP4AB:::ind::D||
Dimethicone_410|ok||||
Choline_salicylate|ok_nutra|PCY1B:::pro::D;ACES:::pro::D;PCY1A:::pro::D;PLD2:::pro::D;CHLE:::pro::D;PLD1:::pro::D;PHOP1:::pro::D;ACHA7|CEPT1:::sub::D;CHKB:::sub::D;CLAT:::sub::D;CHKA:::sub::D;CHDH:::sub::D|S22A2:::inh::D;S22A1:::inh::D;S22A3:::inh::D;S22A5:::inh::D;S22A4:::inh::D;CTL1:::sub::D;CTL4:::sub::D;CTL2:::sub::D;CTL3:::sub::D;SC5A7:::sub::D|
Pentetic_acid|ok|Transuranium_elements:::chel::D|||A1AT:::sub::D
Burosumab|ok_inv|Fibroblast_growth_factor_23:::ant::D|||
Sodium_bisulfite|ok||||
Ox_bile_extract|ok_exp_inv||||
Bromotheophylline|ok||CP1A2:::sub::D||
Fosnetupitant|ok|NK1R:::ant::D|CP3A4:::inh::D||
Benzoin|ok_exp||||
Typhoid_vaccine|ok||||
Nordazepam|exp||||
Acetyl_sulfisoxazole|ok_vet|DHPS::ECOLI:inh::D|CP2C9:::inh::D||
Erenumab|ok_inv|CALRL|||
Fremanezumab|ok_inv|CALCA:::abo::D;CALCB:::abo::D|||
Galcanezumab|ok_inv|CALCA:::abo::D;CALCB:::abo::D|||
Dichlorobenzene|ok_exp||CP2E1:::sub::D||
Sodium_zirconium_cyclosilicate|ok_inv||||
Imidurea|ok_exp||||
Medronic_acid|ok_inv||||
Betiatide|ok_exp||||
Bisphenol_A_diglycidyl_ether|ok_exp||||
Butylparaben|ok_exp||||
Cianidanol|ok_out||||
Dimercaptosuccinic_acid|ok_exp||||
1_2_icosapentoyl_sn_glycero_3_phosphoserine|ok_exp||||
1_2_Distearoyllecithin|ok_exp||||
Pork_Collagen|ok_inv||||
Soy_isoflavones|ok_exp||||
Linoleic_acid|ok_exp||||
Sodium_1_2_Dipalmitoyl_sn_glycero_3_phospho_1_rac_glycerol|ok_exp||||
Tetrakis_2_methoxyisobutylisocyanide_copper_I_tetrafluoroborate|ok||||
alpha_Arbutin|ok_exp||||
Butylene_glycol|ok_exp||||
Human_vaccinia_virus_immune_globulin|ok||||
Black_widow_spider_antivenin_equine|ok||||
Viper_antivenom|ok||||
Human_botulinum_neurotoxin_A_B_immune_globulin|ok||||
Silodrate|ok_exp||||
Phenylethyl_resorcinol|ok_exp||||
Racementhol|ok_exp||||
Hydroxyethyl_ethylcellulose|ok_exp||||
p_Phenylenediamine|ok_exp||||
Distearyldimonium|ok_exp||||
Human_albumin_microspheres|ok_exp||||
Chloric_acid|ok_exp||||
Phosphorus|ok_exp||||
Synthetic_camphor|ok_exp||||
Microcrystalline_cellulose|ok_exp_inv||||
Oxidronic_acid|ok||||
Northern_bluefin_tuna|ok||||
Anthoxanthum_odoratum|ok||||
Betula_lenta_whole|ok||||
Culex_pipiens|ok||||
Rumex_acetosella_whole|ok||||
Rumex_crispus_top|ok||||
Sarocladium_strictum|ok||||
Salix_nigra_bark|ok||||
Artemisia_vulgaris_root|ok_inv||||
Penicillium_glaucum|ok||||
Evernia_prunastri|ok||||
Diazolidinylurea|ok_exp||||
Dipentamethylenethiuram_disulfide|ok_exp||||
alpha_Amyl_cinnamaldehyde|ok_exp||||
Benzylparaben|ok_exp||||
Propylparaben|ok_exp||||
Tetramethylthiuram_monosulfide|ok_exp||||
Phleum_pratense_top|ok||||
Nickel_sulfate|ok_exp||||
Lanolin_alcohols|ok_exp||||
Dichromate|ok_inv||||
Geraniol|ok_exp||||
Cinnamaldehyde|ok_exp||||
Aripiprazole_lauroxil|ok_inv|DRD2:::pag::D;5HT1A:::pag::D;5HT2A:::ant::D;5HT1B;5HT1D;5HT1E;DRD1;DRD5;DRD3;DRD4;5HT2C;5HT3A;5HT6R;5HT7R;HRH1:::ant::D;ADA1A:::ant::D;ADA1B:::ant::D;ADA2A;ADA2B;ADA2C;ACM1;ACM2;ACM3;ACM4;ACM5|CP3A4:::sub::D;CP2D6:::sub::D;CP3A5:::sub::D;CP3A7:::sub::D||ALBU:::bin::D
Cinnamyl_alcohol|ok_exp||||
Hydroxycitronellal|ok_exp||||
Isoeugenol|ok_exp||||
Ethylenediamine|ok_exp||||
P_Tert_Butylphenol_Formaldehyde_Resin_Low_Molecular_Weight|ok_exp||||
Diphenylguanidine|ok_exp||||
N_N_diphenyl_1_4_phenylenediamine|ok_exp||||
Ditiocarb_Zinc|ok_exp||||
Zinc_Dibutyldithiocarbamate|ok_exp||||
4_Isopropylamino_diphenylamine|ok_exp||||
N_Cyclohexyl_N_phenyl_1_4_phenylenediamine|ok||||
Methylchloroisothiazolinone|ok_exp||||
Quaternium_15|ok_exp||||
Bromothalonil|ok_exp||||
Thiohexam|ok_exp||||
2_2_Dibenzothiazyl_disulfide|ok_exp||||
Morpholinylmercaptobenzothiazole|ok_exp||||
Disperse_Blue_106|ok_exp||||
Cobalt_chloride|ok_exp||||
Fanolesomab|ok_exp||||
Methylparaben|ok||||
Telotristat|exp||||
Bifidobacterium_longum_infantis|ok_exp||||
Albumin_Aggregated|ok||||
Quinoline_Yellow_WS|ok_exp||||
Egg_phospholipids|ok_exp_inv||||
Bilberry|ok_exp||||
Echinacea_angustifolia_root|ok_exp||||
Echinacea_purpurea_flowering_top|ok_exp||||
Echinacea_purpurea|ok_exp||||
Echinacea|ok_exp||CP3A4:::ind::D||
Caviar_unspecified|ok_exp||||
Honey|ok_exp||||
Snail_unspecified|ok_exp||||
Jojoba_oil|ok_exp_inv||||
Avena_sativa_flowering_top|ok_exp||||
Aloe_vera_flower|ok_exp||||
Centella_asiatica|ok_exp_inv||||
Aloe_ferox_leaf|ok_exp||||
Elm|ok_exp||||
Bird_pepper|ok_exp||||
Calendula_officinalis_flower|ok_exp||||
Rumex_crispus_whole|ok_exp||||
Ocimum_tenuiflorum_top|ok_exp||||
Salix_alba_bark|ok_exp||||
Indian_frankincense|ok_exp_inv||||
Turmeric|ok_exp_inv||||
Carthamus_tinctorius_flower_bud|ok_exp||||
Corydalis_ambigua_tuber|ok_exp||||
Lonicera_caprifolium_flower|ok_exp||||
Angelica_archangelica_root|ok_exp||||
Kaempferia_galanga_root|ok_exp||||
Larix_sibirica_wood|ok_exp||||
Wormwood|ok_exp||||
Eleuthero|ok_exp||||
Glycyrrhiza_glabra|ok_exp||||
Eucalyptus_globulus_leaf|ok_exp||||
Apricot_kernel_oil|ok_exp||||
Purslane|ok_exp||||
Heterotheca_inuloides_flower|ok_exp||||
Inonotus_obliquus_fruiting_body|ok_exp||||
Nelumbo_nucifera_flower|ok_exp||||
Atractylodes_lancea_root_oil|ok_exp||||
Scutellaria_lateriflora|ok_exp||||
Arnica_montana_flower|ok_exp||||
Equisetum_arvense_top|ok_exp||||
Inula_helenium_root|ok_exp||||
Usnea_barbata|ok_exp||||
Azadirachta_indica_leaf|ok_exp||||
Zanthoxylum_clava_herculis_whole|ok_exp||||
Chamomile|ok_exp_inv||||
Saw_palmetto|ok_exp_inv||||
Rice_bran|ok_exp||||
Milk_thistle|ok_exp_inv||||
Influenza_A_virus_A_California_7_2009_H1N1_like_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_179A_H1N1_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Victoria_210_2009_X_187_H3N2_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Brisbane_60_2008_hemagglutinin_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_A_virus_A_Victoria_361_2011_IVR_165_H3N2_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Texas_6_2011_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Bordetella_pertussis_toxoid_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_X_223A_H3N2_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Christchurch_16_2010_NIB_74_H1N1_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_X_223_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_H1N1_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Victoria_361_2011_H3N2_live_attenuated_antigen|ok||||
Influenza_B_virus_B_Wisconsin_1_2010_live_attenuated_antigen|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_BX_51B_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Brisbane_10_2010_H1N1_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_X_223A_H3N2_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_BX_51B_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Switzerland_9715293_2013_NIB_88_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_181_H1N1_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Switzerland_9715293_2013_NIB_88_H3N2_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Brisbane_9_2014_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_South_Australia_55_2014_IVR_175_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Human_adenovirus_e_serotype_4_strain_cl_68578_antigen|ok||||
Human_adenovirus_b_serotype_7|ok||||
Influenza_A_virus_A_Victoria_361_2011_IVR_165_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Hubei_Wujiagang_158_2009_BX_39_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_X_263B_H3N2_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_179A_H1N1_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Switzerland_9715293_2013_NIB_88_H3N2_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_H3N2_recombinant_hemagglutinin_antigen|ok||||
Influenza_B_virus_B_Brisbane_60_2008_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Christchurch_16_2010_NIB_74XP_H1N1_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_South_Australia_55_2014_H3N2_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Utah_9_2014_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Michigan_45_2015_X_275_H1N1_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Michigan_45_2015_H1N1_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_X_263B_H3N2_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Slovenia_2903_2015_H1N1_live_attenuated_antigen|ok||||
Influenza_A_virus_A_New_caledonia_71_2014_H3N2_live_attenuated_antigen|ok||||
Neisseria_meningitidis_group_a_capsular_oligosaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Neisseria_meningitidis_group_c_capsular_oligosaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Neisseria_meningitidis_group_w_135_capsular_oligosaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Neisseria_meningitidis_group_y_capsular_oligosaccharide_diphtheria_crm197_protein_conjugate_antigen|ok||||
Influenza_A_virus_A_Singapore_gp1908_2015_IVR_180_H1N1_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_gp1908_2015_IVR_180_H1N1_hemagglutinin_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Singapore_gp1908_2015_IVR_180_H1N1_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_gp2050_2015_H3N2_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Hong_Kong_259_2010_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_H3N2_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_gp1908_2015_IVR_180_H1N1_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_X_263B_H3N2_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Brisbane_60_2008_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Singapore_GP1908_2015_IVR_180A_H1N1_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Brisbane_46_2015_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_BVR_1B_hemagglutinin_antigen_propiolactone_inactivated|ok||||
Vibrio_cholerae_CVD_103_HgR_strain_live_antigen|ok_inv||||
Influenza_A_virus_A_California_7_2009_H1N1_like_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Victoria_210_2009_X_187_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_South_Dakota_6_2007_H1N1_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Uruguay_716_2007_H3N2_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Perth_16_2009_H3N2_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Victoria_361_2011_IVR_165_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Texas_6_2011_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_X_223A_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_BX_51B_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_181_H1N1_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Brisbane_9_2014_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_X_263B_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Michigan_45_2015_X_275_H1N1_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_X_263B_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_gp1908_2015_IVR_180_H1N1_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_gp1908_2015_IVR_180_H1N1_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Singapore_GP1908_2015_IVR_180_H1N1_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_GP2050_2015_H3N2_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Hong_Kong_259_2010_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_H3N2_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_GP1908_2015_IVR_180_H1N1_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Hong_Kong_4801_2014_X_263B_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Singapore_GP1908_2015_IVR_180A_H1N1_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Brisbane_46_2015_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Phuket_3073_2013_BVR_1B_antigen_propiolactone_inactivated|ok||||
Beroctocog_alfa|ok_inv||||
DL_alpha_Tocopherol|ok_exp_inv||||
DL_alpha_tocopheryl_acetate|ok_exp||||
Povidone_K30|ok_exp||||
Calcium_phosphate_dihydrate|ok|CASR;CALR;CIB1;PDCD6;SORCN;CHP1;SPRC;CALX;FBN2;S100B;CASQ2;RGN;PEF1;S10A6;TCTP;CIB2;S10AD;CASQ1;NUCB1;NUCB2;CALM1;FBN3;GRAN;CAPS1;CALM2;CALM3;S10AG;CALB2;CAYP1;CAPS2;CALR3;NRX1A;NCS1||S20A1;S20A2;NPT2A;NPT2B;NPT2C;TRPV6;NAC1;TRPV5;RYR1;RYR2;PK2L1;RYR3;PK1L3;CTSR1;CAC1C;CAC1A;CAC1G;CAC1E|CALB1;S100G;ALBU
Sodium_ascorbate|ok_nutra||||
Calcium_ascorbate|ok_nutra||||
Magnesium_ascorbate|ok_nutra||||
Zinc_ascorbate|ok_nutra||||
Niacinamide_ascorbate|ok_nutra||||
Zinc_acetate|ok_inv|BKRB1;MGMT;ALDOA;EF1A1;ENOA;G3PT;NDKA;PDIA1;PDIA3;PRDX1;SERB;TPIS;EFTU;ESR1;IL3;MT2;CCS;HDAC1;HDAC4;3MG;SEMG1;SODC;HDAC8;SIVA;GLRA1;MDM2;INS;UTRO;ACY2;S10A8;S10A9;MMP9;P73;S10A2;P53;MT3;PDCD6;DAND5;MT1A;A1BG;A2MG;ANGT;FETUA;SAMP;APOA1;APOA2;APOA4;APOBR;APOE;APOL1;C1QB;C1QC;C1R;C1S;CO3;CO4B;C4BPA;C4BPB;CO5;BRCC3;CO8A;CO8B;CO8G;CFAB;CFAH;CFAI;CLUS;CERU;CBPN;CPN2;DCD;DESP;FA12;F13B;THRB;FCN3;FIBA;FINC;GELS;HBA;HBB;HPTR;HORN;ALS;IGHA1;IGHM;KV117;KV320;LV321;ITIH1;ITIH2;ITIH3;ITIH4;IGJ;PLAK;KLKB1;KNG1;K2C1;K1C10;K1C14;K1C16;K22E;K2C5;K2C6A;K1C9;A1AG2;PGRP2;PON1;PZP;S10A7;SEPP1;A1AT;AACT;KAIN;CBG;HEP2;SHBG;TRFE;TTHY;VTNC;APLP1;APLP2;A4;PARP1|CAH1:::lig::D;CBPE:::inh::D;ADH1G:::lig::D;IDE:::lig::D;SODC:::lig::D||
Ferrous_gluconate|ok|TFR1;EGLN1;HDAC8;AHSP;HBA;FRDA;FRIH;FEN1;NEIL1;NEIL2;DPOLB;CERU;TRFE|||
Ferrous_succinate|ok|TFR1;EGLN1;HDAC8;AHSP;HBA;FRDA;FRIH;FEN1;NEIL1;NEIL2;DPOLB;CERU;TRFE|||
Ferrous_ascorbate|ok|TFR1;EGLN1;HDAC8;AHSP;HBA;FRDA;FRIH;FEN1;NEIL1;NEIL2;DPOLB;CERU;TRFE|||
Ferrous_fumarate|ok|TFR1;EGLN1;HDAC8;AHSP;HBA;FRDA;FRIH;FEN1;NEIL1;NEIL2;DPOLB;CERU;TRFE|||
Sodium_molybdate|ok_exp||||
Potassium_acetate|ok_inv|AT1A1|||
Potassium_sulfate|ok_inv|AT1A1|||
Potassium|ok_exp|AT1A1:::reg::D||AT1A1:::sub::D;S12A1:::lig::D|
Ferrous_glycine_sulfate|ok|TFR1;EGLN1;HDAC8;AHSP;HBA;FRDA;FRIH;FEN1;NEIL1;NEIL2;DPOLB;CERU;TRFE|||
Sodium_phosphate_dibasic|ok|||S20A1;S20A2;NPT2A;NPT2B;NPT2C|
Sodium_phosphate_monobasic_unspecified_form|ok|||S20A1;S20A2;NPT2A;NPT2B;NPT2C|
Sodium_phosphate_dibasic_unspecified_form|ok_exp||||
Sodium_borate|ok_exp||||
Lithium_hydroxide|ok_out||||
Lithium_citrate|ok|IMPA2;IMPA1;GSK3B;GRIA3|||
Lithium_succinate|exp|IMPA2;IMPA1;GSK3B;GRIA3|||
Lithium_carbonate|ok|IMPA2;IMPA1;GSK3B;GRIA3||SCNNA;SCNNB;SCNNG|
Mometasone_furoate|ok_inv_vet|GCR;PRGR|CP2C8:::inh::D;CP3A4:::sub_ind::D;CP3A5:::ind::D||
Magnesium|ok_exp_inv||||ALBU
Magnesium_levulinate|nutra|AT1A1|||
Magnesium_lactate|nutra|AT1A1|||
Aluminium_phosphate|ok_inv|TRFE;AT1A1;KLK1;A4|||ALBU
Aluminum_acetate|ok_inv|TRFE;AT1A1;KLK1;A4|||ALBU
Tetraferric_tricitrate_decahydrate|ok|FHUD::ECOLI:::D;TFR1|||TRFE;ITB3;CALR
Chromic_nitrate|ok|CYB5|||TRFE
Chromium_gluconate|ok|CYB5|||TRFE
Chromium_nicotinate|ok_exp|CYB5|||TRFE
Chromous_sulfate|ok|CYB5|||TRFE
Zinc_chloride|ok_inv|BKRB1;MGMT;ALDOA;EF1A1;ENOA;G3PT;NDKA;PDIA1;PDIA3;PRDX1;SERB;TPIS;EFTU;ESR1;IL3;MT2;CCS;HDAC1;HDAC4;3MG;SEMG1;SODC;HDAC8;SIVA;GLRA1;MDM2;INS;UTRO;ACY2;S10A8;S10A9;MMP9;P73;S10A2;P53;MT3;PDCD6;DAND5;MT1A;A1BG;A2MG;ANGT;FETUA;SAMP;APOA1;APOA2;APOA4;APOBR;APOE;APOL1;C1QB;C1QC;C1R;C1S;CO3;CO4B;C4BPA;C4BPB;CO5;BRCC3;CO8A;CO8B;CO8G;CFAB;CFAH;CFAI;CLUS;CERU;CBPN;CPN2;DCD;DESP;FA12;F13B;THRB;FCN3;FIBA;FINC;GELS;HBA;HBB;HPTR;HORN;ALS;IGHA1;IGHM;KV117;KV320;LV321;ITIH1;ITIH2;ITIH3;ITIH4;IGJ;PLAK;KLKB1;KNG1;K2C1;K1C10;K1C14;K1C16;K22E;K2C5;K2C6A;K1C9;A1AG2;PGRP2;PON1;PZP;S10A7;SEPP1;A1AT;AACT;KAIN;CBG;HEP2;SHBG;TRFE;TTHY;VTNC;APLP1;APLP2;A4;PARP1|CBPE:::inh::D;ADH1G:::lig::D;IDE:::lig::D;SODC:::cof::D;CAH2:::cof::D||
Hydrocortisone_aceponate|exp_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub_ind::D;CP3A5:::sub::D;CP3A7:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_acetate|ok_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub_ind::D;CP3A5:::sub::D;CP3A7:::sub::D;C11B1:::sub::D;C11B2:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_butyrate|ok_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub_ind::D;CP3A5:::sub::D;CP3A7:::sub::D;C11B1:::sub::D;C11B2:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_cypionate|ok_inv_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub::D;CP3A5:::sub::D;CP3A7:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_phosphate|ok_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub::D;CP3A5:::sub::D;CP3A7:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_probutate|ok_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub_ind::D;CP3A5:::sub::D;CP3A7:::sub::D;C11B1:::sub::D;C11B2:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_valerate|ok_vet|ANXA1;GCR;DHI2;3BHS1|CP3A4:::sub_ind::D;CP3A5:::sub::D;CP3A7:::sub::D;C11B1:::sub::D;C11B2:::sub::D;CP2C8:::ind::D|MDR1;SO1A2;ABCG2;S22A8|SHBG;CBG
Hydrocortisone_succinate|ok||CP3A4:::sub_ind::D;CP2C8:::ind::D;C11B1:::sub::D;C11B2:::sub::D||
Zinc_sulfate_unspecified_form|ok_exp||||
Gallium_chloride_Ga_67|ok_exp||||
Dotatate|ok_exp||||
Ursadiol|ok_exp||||
Influenza_A_virus_A_Singapore_INFIMH_16_0019_2016_NIB_104_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Maryland_15_2016_BX_69A_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Singapore_INFIMH_16_0019_2016_IVR_186_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Maryland_15_2016_BX_69A_antigen_UV_formaldehyde_inactivated|ok||||
Andexanet_alfa|ok_inv|TFPI1:::inh::D|||
Lavender_oil|ok_exp||||
Brown_iron_oxide|ok_exp||||
Ivosidenib|ok_inv|IDHC:::inh::D|CP3A4:::sub_ind::D;CP2B6:::ind::D;CP2C9:::ind::D;CP2C8:::ind::D|S22A8:::inh::D;MDR1:::inh::D|
Tedizolid|ok_inv||||
Hydroxyprogesterone|exp||CP3A4:::sub::D||
Cobalt|ok_exp||||
Eslicarbazepine|ok|P2RX4|UD11:::sub::D;CP2CJ:::inh::D;CP3A4:::ind::D||
Patisiran|ok_inv|Transthyretin_mRNA:::sup::D|||ALBU:::lig::D;A1AG1:::lig::D
Segesterone_acetate|ok_exp_inv|PRGR:::ago::D;ANDR:::ago::D;GCR:::ago::D|CP3A4:::sub::D||
Plantago_ovata_seed|ok_exp_inv||||
Citrus_bioflavonoids|ok_exp||||
Influenza_A_virus_A_Singapore_INFIMH_16_0019_2016_IVR_186_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Maryland_15_2016_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Singapore_INFIMH_16_0019_2016_IVR_186_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Maryland_15_2016_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Singapore_INFIMH_16_0019_2016_H3N2_recombinant_hemagglutinin_antigen|ok||||
Influenza_B_virus_B_Maryland_15_2016_recombinant_hemagglutinin_antigen|ok||||
Loteprednol|ok_exp||||
Lanadelumab|ok_inv|KLKB1:::inh::D|||
Edetate_calcium_disodium_anhydrous|ok||||
Edetate_disodium_anhydrous|ok_vet|Lead;Iron;Manganese_cation|ADA:::inh::D;PON3:::inh::D;CP19A:::inh::D;CP3A4:::inh::D;PON1:::inh::D||
Barley_malt_syrup|ok||||
Influenza_A_virus_A_Victoria_361_2011_IVR_165_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Hubei_Wujiagang_158_2009_BX_39_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_X_223A_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_BX_51B_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Texas_50_2012_H3N2_live_attenuated_antigen|ok||||
Influenza_B_virus_B_Massachusetts_2_2012_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Victoria_361_2011_IVR_165_H3N2_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Wisconsin_1_2010_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Hubei_Wujiagang_158_2009_BX_39_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Victoria_210_2009_X_187_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_California_7_2009_X_181_H1N1_antigen_UV_formaldehyde_inactivated|ok||||
Serum_horse|ok||||
Influenza_A_virus_A_Victoria_210_2009_X_187_H3N2_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Uruguay_716_2007_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Brisbane_59_2007_H1N1_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Uruguay_716_2007_H3N2_hemagglutinin_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_A_virus_A_Brisbane_59_2007_H1N1_hemagglutinin_antigen_formaldehyde_inactivated|ok_inv||||
Influenza_A_virus_A_Uruguay_716_2007_H3N2_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Brisbane_59_2007_H1N1_antigen_propiolactone_inactivated|ok||||
Oxyphenisatin_acetate|ok_out||||
Prednisolone_phosphate|ok_vet||CP3A4:::ind::D;CP3A5:::ind::D||
Prednisolone_tebutate|ok_vet||||
Diloxanide_furoate|ok||||
Lypressin|ok|V1AR;V2R;V1BR||MRP2|
Methylprednisolone_aceponate|ok_vet||||
Methylprednisolone_hemisuccinate|ok||CP3A4:::ind::D;CP3A5:::ind::D||
Prednisone_acetate|ok_exp_inv||CP3A4:::ind::D;CP3A5:::ind::D||
Dexamethasone_acetate|ok_inv_vet||||
Menadiol_diphosphate|ok_nutra||||
Drostanolone_propionate|ok_ill||||
Chlorphenesin_carbamate|ok_vet_out||||
Paramethasone_acetate|ok||||
Chloramphenicol_palmitate|ok_vet||||
Loperamide_oxide|exp||||
Betamethasone_phosphate|ok_vet||CP3A4:::ind::D;CP3A5:::ind::D||
Estramustine_phosphate|ok_inv||||
Gestonorone_caproate|ok||||
Cortisone|exp||CP3A4:::ind::D;CP3A5:::ind::D||
Calcium_polycarbophil|ok||||
Adenovirus_type_7_vaccine_live|ok||||
Rosemary_oil|ok_exp||||
Ginger_oil|ok_exp||||
Willow_bark|ok_exp||||
Turmeric_oil|ok_exp||||
Atractylodes_lancea_root|ok_exp||||
Beef_liver|ok_exp||||
Ferric_oxyhydroxide|ok_exp||||
Influenza_A_virus_A_Singapore_INFIMH_16_0019_2016_H3N2_live_attenuated_antigen|ok||||
Influenza_B_virus_B_Colorado_06_2017_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Brisbane_59_2007_H1N1_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Uruguay_716_2007_H3N2_hemagglutinin_antigen_UV_formaldehyde_inactivated|ok||||
Damoctocog_alfa_pegol|ok_inv|FA8:::bin::D|||
Sodium_metavanadate|ok_exp||||
Dexamethasone_metasulfobenzoate|ok_exp||||
Cemiplimab|ok_inv|PDCD1:::inh::D|||
Tosylchloramide|exp||||
Bean|ok||||
Camponotus_pennsylvanicus|ok||||
Vaccinia_virus_strain_new_york_city_board_of_health_live_antigen|ok||||
Elapegademase|ok||||
Inotersen|ok_inv|Transthyretin_mRNA:::inh::D|||
Bentazepam|exp||||
Larotrectinib|ok_inv|NTRK1:::inh::D;NTRK2:::inh::D;NTRK3:::inh::D|CP3A4:::sub::D||
Emapalumab|ok_inv|IFNG:::neu::D|||
Cefamandole_nafate|ok||||
Calaspargase_pegol|ok|L_asparagine:::degr::D|||
Tagraxofusp|ok_inv|IL3RA:::bin::D;ARL2:::bin::D|||
Ceftobiprole_medocaril|exp_inv||||
Turoctocog_alfa_pegol|ok|FA9:::act::D;FA10:::act::D;THRB:::bin::D|PROC:::sub::D;FA10:::sub::D||VWF:::bin::D
Hyaluronidase|ok||||
Luteinizing_hormone|ok||||
Polymyxin_B|ok_vet|Bacterial_outer_membrane::Bacteria:destbz::D||S15A2|
Polygala_senega_root|exp||||
Mecasermin_rinfabate|ok|IGF1R:::ago::D;INSR;MPRI|||
Racephedrine|ok_exp||||
Hydroxystilbamidine|ok|DNA|||
Solriamfetol|ok|SC6A3;SC6A2||S22A2;S22A4;S22A5|
Agrostis_gigantea_top|ok||||
Catfish|ok||||
Red_pepper|ok||||
Risankizumab|ok_inv|IL12B:::inh::D|||
Cycloguanil|ok||||
Dengue_tetravalent_vaccine_live|ok||||
Diroximel_fumarate|ok_inv|ACH10:::ago::D|Liver_esterases:::sub::D||
Brolucizumab|ok_inv|VEGFA:::inh::D|||
Cefiderocol|ok_inv|Cell_division_protein::PSEAI:inh::D;PBPA::PSEAE:inh::D;Penicillin_binding_protein_1B::PSEAI:inh::D;Penicillin_binding_protein_2::PSEAI:inh::D;DACB::ECOLI:inh::D||MEXA::PSEAE:sub::D;FIU::ECOLI:sub::D;CIRA::ECOLI:sub::D;A0A0H2ZGX7:::sub::D|ALBU:::lig::D
Bermekimab|inv||||
Etirinotecan_pegol|inv||||
Trastuzumab_deruxtecan|ok_inv|FCGR1:::abo::D;TOP1:::inh::D|LYAG:::sub::D;TOP1:::inh::D;CATB:::sub::D;CATL1:::sub::D;CP3A4:::sub::D|MDR1:::sub::D;SO1B1;SO1B3:::sub::D;S47A2:::sub::D;MRP1:::sub::D;ABCG2:::sub::D|
Voxelotor|ok_inv|HBA:::bin::D|CP3A4:::sub::D;CP2C9:::sub::D;CP2B6:::sub::D;CP2CJ:::sub::D||
Zanubrutinib|ok_inv|BTK:::inh::D;EGFR:::inh::D;ERBB2:::inh::D;ERBB4:::inh::D;ITK:::inh::D;BMX:::inh::D;JAK2:::inh::D;TEC:::inh::D;BLK:::inh::D;JAK3:::inh::D;PTK6:::inh::D;FGR:::inh::D;FRK:::inh::D;LCK:::inh::D;TXK:::inh::D|CP3A4:::sub::D;CP2B6:::ind::D|MDR1:::sub::D|
Givosiran|ok_inv|ALAS1_mRNA:::cli::D|||
Upadacitinib|ok_inv|JAK1:::inh::D|CP3A4:::sub::D;CP2D6:::sub::D|MDR1:::inh::D;ABCG2:::inh::D;SO1B1:::inh::D|
Ropeginterferon_alfa_2b|inv||CP1A2:::inh::D||
Thyrotropin|inv||||
Crizanlizumab|ok_inv|LYAM3:::inh::D|||
Pertussis_vaccine|ok_inv||||
Pegteograstim|inv||||
Hydroquinidine|inv||||
Ubrogepant|ok_inv|CALRL:::ant::D|CP3A4:::sub::D;CP2C8:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D;AOFA:::inh::D;UD11:::inh::D;CP2D6:::inh::D|MDR1:::sub::D;ABCG2:::sub::D;SO1B1:::inh::D;SO1B3:::inh::D;S22A6:::sub::D;S22A2:::inh::D|
Elexacaftor|ok_inv|CFTR:::mod::D|CP3A4:::inh::D;CP3A5:::sub::D;CP1A2:::inh::D;CP2B6:::inh::D;CP2C8:::inh::D;CP2C9:::inh::D;CP2CJ:::inh::D;CP2D6:::inh::D|SO1B1:::inh::D;SO1B3:::inh::D;MDR1:::inh::D|ALBU:::sub::D
Benzhydrocodone|ok||||
Cinoxate|ok||||
Haemagglutinin_strain_B_Victoria|ok||||
Haemagglutinin_strain_B_Yamagata|ok||||
Haemagglutinin_strain_A_H3N2|ok||||
Haemagglutinin_strain_A_H1N1|ok||||
Alloin|ok_exp||||
Frangula_purshiana_bark|ok_exp||||
Zirconium_chloride_hydroxide|ok_exp||||
Resorcinol_monoacetate|ok_exp||||
Fish_liver_oil|ok_exp||||
Haemagglutinin_strain_B|ok||||
Modified_vaccinia_ankara|ok||||
VIBRIO_CHOLERAE_INABA_6973_E1_TOR_BIOTYPE_FORMALIN_INACTIVATED|ok||||
VIBRIO_CHOLERAE_INABA_48_CLASSICAL_BIOTYPE_HEAT_INACTIVATED|ok||||
VIBRIO_CHOLERAE_OGAWA_50_CLASSICAL_BIOTYPE_HEAT_INACTIVATED|ok||||
VIBRIO_CHOLERAE_OGAWA_50_CLASSICAL_BIOTYPE_FORMALIN_INACTIVATED|ok||||
Edotreotide_gallium_Ga_68|ok|SSR2:::lig::D;SSR5:::lig::D;SSR3:::lig::D;SSR1:::lig::D|||
Smallpox_and_Monkeypox_Vaccine_Live_Non_replicating|ok||||
Influenza_A_virus_A_Brisbane_02_2018_IVR_190_H1N1_antigen_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Kansas_14_2017_X_327_H3N2_antigen_propiolactone_inactivated|ok||||
Baccharis_sarothroides_whole|ok||||
Amaranthus_hybridus_pollen|ok||||
Acacia_dealbata_pollen|ok||||
Influenza_A_virus_A_Idaho_07_2018_H1N1_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_A_virus_A_Indiana_08_2018_H3N2_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Singapore_INFTT_16_0610_2016_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Iowa_06_2017_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Alnus_serrulata_pollen|ok||||
Prosopis_velutina_seed|ok||||
Gibberella_fujikuroi|ok||||
Mucor_circinelloides_f_circinelloides|ok||||
Influenza_A_virus_A_Switzerland_3330_2017_H1N1_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Kansas_14_2017_H3N2_live_attenuated_antigen|ok||||
Influenza_A_virus_A_Brisbane_02_2018_IVR_190_H1N1_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Kansas_14_2017_X_327_H3N2_antigen_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Brisbane_02_2018_H1N1_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Kansas_14_2017_H3N2_recombinant_hemagglutinin_antigen|ok||||
Influenza_A_virus_A_Brisbane_02_2018_IVR_190_H1N1_antigen_UV_formaldehyde_inactivated|ok||||
Influenza_A_virus_A_Kansas_14_2017_X_327_H3N2_antigen_UV_formaldehyde_inactivated|ok||||
Cyd_dengue_virus_serotype_1_live_attenuated_antigen|ok||||
Cyd_dengue_virus_serotype_2_live_attenuated_antigen|ok||||
Cyd_dengue_virus_serotype_3_live_attenuated_antigen|ok||||
Cyd_dengue_virus_serotype_4_live_attenuated_antigen|ok||||
Mucor_circinelloides_f_lusitanicus|ok||||
Eurotium_amstelodami|ok||||
Onasemnogene_abeparvovec|ok||||
Leucanthemum_vulgare_pollen|ok||||
Trifolium_pratense_pollen|ok||||
Colchiceine|ok_exp||||
Eucalyptus_gum|ok_exp||||
Sea_scallop|ok||||
Northern_brown_shrimp|ok||||
Rainbow_trout|ok||||
Yellowfin_tuna|ok||||
Atlantic_mackerel|ok||||
Pacific_ocean_perch|ok||||
Myristica_fragrans_fruit|ok||||
Pisum_sativum_whole|ok||||
Skim_milk|ok||||
Black_sea_bass|ok||||
Channel_catfish|ok||||
Atlantic_halibut|ok||||
Influenza_A_virus_A_North_carolina_04_2016_H3N2_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Iowa_06_2017_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Influenza_B_virus_B_Singapore_INFTT_16_0610_2016_hemagglutinin_antigen_MDCK_cell_derived_propiolactone_inactivated|ok||||
Prednisolone_acetate|ok_vet|GCR:::ago::D|CP3A4:::sub_ind::D|SO1A2:::inh::D;MDR1:::sub::D|CBG:::bin::D;ALBU:::bin::D
Padeliporfin|exp||||
Ethyl_salicylate|ok_exp||||
Desfesoterodine|exp||||
Cucurbita_pepo_subsp_ovifera_whole|ok||||
Golodirsen|ok|DMD:::ind::D|||
Brilliant_blue_G|ok|Internal_limiting_membrane_ILM:::bin::D|||
Ebola_Zaire_vaccine_live_attenuated|ok||||
Ferric_maltol|ok||||
