name|status|tar|enz|tra|car
Drug1|ok|TAR1:::inh:<9.5:D;TAR2:::inh:<7.0:D;TAR3:::inh:<10:D;TAR4:::inh:8:D;TAR5:::inh:8:D;TAR6:::inh:7:D;TAR7:::inh:8:D;TAR8:::inh:<6:D;TAR9:::inh:9:D;TAR10:::inh:<9:D;TAR11:::inh:>7:D;TAR12:::inh:>10:D;TAR13:::inh:<8:D;TAR14:::inh:>10:D;TAR15:::inh:>8:D;TAR16:::inh:>7:D;TAR17:::inh:10:D;TAR18:::inh:>10:D;TAR19:::inh:7:D;TAR20:::inh:>9:D;TAR21:::inh::D;TAR22:::inh:<6:D;TAR23:::inh::D|||
Drug2|ok|TAR1:::inh:<7.0:D;TAR2:::inh:<9.5:D;TAR3:::inh:8:D;TAR4:::inh:<10:D;TAR5:::inh:7:D;TAR6:::inh:8:D;TAR7:::inh:<6:D;TAR8:::inh:8:D;TAR9:::inh:9:D;TAR10:::inh:>7:D;TAR11:::inh:<9:D;TAR12:::inh:<8:D;TAR13:::inh:>10:D;TAR14:::inh:>8:D;TAR15:::inh:>10:D;TAR16:::inh:10:D;TAR17:::inh:>7:D;TAR18:::inh:7:D;TAR19:::inh:>10:D;TAR20:::inh::D;TAR21:::inh:>9:D;TAR22:::inh::D;TAR23:::inh:<6:D|||
